module green_reverse(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100011111010011101100101010101010010110101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011011010001010101110111011001111001011110001,
	240'b111100001110101011000101110010011110001111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100001101110111000001110001011110111111110000,
	240'b111011111011110111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101100100011110000,
	240'b110000111100111011111111111101111011110110100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100001100111101001111010100001101000111100101011111110111111101100001011000011,
	240'b100111101111000111111110100111110101000101001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111101011000011110110111100101010111010011100101011110111110111111111101111110011011,
	240'b101011011111111111101011011000110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101111110011001100101010100100100111101111110111111001110111110110011,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110010111010011111111110111001010101100101000001110011111101101111000010111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000100110101101110011111111101010100101000101110010111101101111000010111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110110110001011110011100011111111011000010101101110111101101111000010111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111011111011110110101111011111010110101101101111101101111000010111110,
	240'b101101001111111111011111010111100101001101010011010100000100111101001111010100000101000101010011010101000101010101010101010101010101010101010101010101010101010101010010100001111111011111101110101101101000010001110000111101101111000010111110,
	240'b101101001111111111011111010111100101000001011110100010001001110110011010100100010111110001100110010101110101000001010010010101010101010101010101010101010101010101010101010100011001100011111011111010011001111101110101111101011111000010111110,
	240'b101101001111111111011111010110100111010111010101111111001111111111111111111111111111100011101100110010101001110101101011010100110101001001010101010101010101010101010101010101000101001010101101111111111100100101110011111101011111000010111110,
	240'b101101001111111111011100011101001110001111111111111111111111111111111111111111111111111111111111111111111111111111101100101101010110110101010001010101000101010101010101010101010101001001111001101101101001000101110011111101011111000010111110,
	240'b101101001111111111011100101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110011010010101110101001001010101010101010101010101010101010100100100111101110011111101101111000010111110,
	240'b101101001111111111101001111011101111111111111111111111111111111111111111111111111111110111111101111111011111110111111011111111111111111111111110101111110110001001010001010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111110001111110011111111111111111111111111111111111111111111110001001110010001000100010101000100111000100111111111111111111111111111111111101010001101001010100010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111110010111110011111111111111111111111111111111111111111111101010110101001001101010011010110011111101010111111111111111111111111111111111111111111010111011010000101000101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111101111111110001111111111111111111111111111111111111111111101010110111001010010010101000101100010110001111111111111111111111111111111111111111111111111110011010101110101010011010101010101000101110011111101101111000010111110,
	240'b101101001111111111101011111101001111111111111111111111111111111111111111111101010110110001001110010101010101001101011000101111011111111111111111111111111111111111111111111111111011000001010011010101000101000101110011111101101111000010111110,
	240'b101101001111111111100101111001011111111111111111111111111111111111111111111100111000010010001100010101000101010001010010010111111100101111111111111111111111111111111111111111111111100110000101010100000101000101110011111101101111000010111110,
	240'b101101001111111111011110110011111111111111111111111111111111111111111111111101111101101111101010100101010101000001010101010100010110010111011000111111111111111111111111111111111111111111011001010111010101000001110011111101101111000010111110,
	240'b101101001111111111011001101011101111111111111111111111111111111111111111111111111101010101111100110110011000100101010000010101010101000101101110111000101111111111111111111111111111111111111111100110010100110001110011111101101111000010111110,
	240'b101101001111111111011010100010001111101011111111111111111111111111111111111111111010011101001010011111111101101101111100010100000101010101010000100000111111100011111111111111111111111111111111110111000101101001110001111101101111000010111110,
	240'b101101001111111111011101011010001110000011111111111111111111111111111111111111111001101101001111010100001000101111010111011100010101000101010100010101111101010111111111111111111111111111111111111111011000011001101110111101101111000010111110,
	240'b101101001111111111011110010110101011000011111111111111111111111111111111111111111010111001001111010101000101000110011001110100110110011101010001010100101011111011111111111111111111111111111111111111111011101001110001111101011111000010111110,
	240'b101101001111111111011111010110100111010111110110111111111111111111111111111111111110000101100010010100100101010001010011101010001100101001011111010100001100011011111111111111111111111111111111111111111110010010000001111101001111000010111110,
	240'b101101001111111111011111010111010101001111000011111111111111111111111111111111111111111110111110010110010101001101010100010101101011011010111101011011011110100111111111111111111111111111111111111111111111100010011101111100011111000010111110,
	240'b101101001111111111011111010111100100111101111000111101011111111111111111111111111111111111111111101011110101010001010100010100110101101010111110111001001110011011111101111111111111111111111111111111111111111110111101111100011111000010111110,
	240'b101101001111111111011111010111100101001101010010101011111111111111111111111111111111111111111111111111011010000101010010010101000101001001100100101000011001101111111110111111111111111111111111111111111111111111011001111100101111000010111110,
	240'b101101001111111111011111010111100101001101010011011000011101101111111111111111111111111111111111111111111111100010010011010100010101010101010100010011011000110111111111111111111111111111111111111111111111111111101010111101001111000010111110,
	240'b101101001111111111011111010111100101001101010101010100010111100011101110111111111111111111111111111111111111111111110011100010000101001101010101010100001000111011111111111111111111111111111111111111111111111111101111111101111110111110111110,
	240'b101101001111111111011111010111100101001101010101010101010101000010001100111101001111111111111111111111111111111111111111110101000101100001001111010011001000101111111111111111111111111111111111111111111111111111110010111110011110111110111110,
	240'b101101001111111111011111010111100101001101010101010101010101010001010001100011111111001011111111111111111111111111111011101010010111011001111000011101001010011011111111111111111111111111111111111111111111111111110010111110011110111110111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010100010100011000001111100110111111111111111111111101111101011111011011110111111101101111100111111111111111111111111111111111111111111111111111101000111101001111000010111110,
	240'b101101001111111111011111010111100100111101010000010101000101010101010101010101010101000101101100110000011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010111100011111000010111110,
	240'b101101001111111111011110011001001001011010100010011010000101001101010101010101010101010101010001010101111000101011010011111111001111111111111111111111111111111111111111111111111111111111111111111111111101001101111110111101001111000010111110,
	240'b101101001111111111011101011010101110100111111110100001010100111101010101010101010101010101010101010101000101000001011100100001111100000111100110111111001111111111111111111111111111111111111111110101100110110101101111111101101111000010111110,
	240'b101101001111111111011101011010101100011011111011111001000110111001010001010101010101010101010101010101010101010101010100010100000101001101100101011111101001100010101100101101101011010010010000010111110100111001110011111101101111000010111110,
	240'b101101001111111111011110011000001001000011000010111111111101100001100110010100110101010101010101010101010101010101010101010101010101010101010011010100010101000001010000010100000101000001010000010100110101000101110011111101101111000010111110,
	240'b101101001111111111011110010111011100111111010100110001101111111110110011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111011110010110111011000111111111110001111101001011001000010101010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111011111010111000110001111010110111111111100010010001110010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111011111010111100100111101101101110111111111110011001001010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101011111111111111100111011000010101001101001111100001001111111111100110010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001111001111110101111000010110110,
	240'b100111101111010011111100100100010100111001001101011000011000110010000001010100100100111101010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110101000110110000111111111110001110011011,
	240'b101110011101010111111111111100001010011010001100100011001000100010001001100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011011011011111010111111111100011010110111,
	240'b111011001011100111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100001011101100,
	240'b111110001110110010111100110101001111000011111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110101011001110110001001111001111111000,
	240'b111111111111111111100101101000001001110010110001101100111011001110110011101100111011001110110011101100101011001010110010101100101011001110110011101100111011001110110011101100111011001010110011101011011001011110110110111110111111111111111111,
	240'b111100011111010011101100101010101010010110101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011011010001010101110111011001111001011110001,
	240'b111100001110101011000101110010011110001111110000111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100001101110111000001110001011110111111110000,
	240'b111011111011110111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101100100011110000,
	240'b110000111100111011111111111110111101111011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110011101100111011010000110100011110010111111111111111101100001011000011,
	240'b100111101111000111111111110011111010100010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101011101111011011110010101011101001101010101111011110111111111101111110011011,
	240'b101011011111111011110101101100011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111110111111001010110010101010001010011110111110111111101110111110110011,
	240'b101101001111111111101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111101001111111111011100101010111010011110111001111110111110111110111110,
	240'b101101001111111111101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000110011011110111011111111110101001010100010111001111110111110111110111110,
	240'b101101001111111111101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111011001101110111110001111111101100001010110111111110111110111110111110,
	240'b101101001111111111101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101100111011101111101111011010111101111101011010110110111110111110111110111110,
	240'b101101001111111111101111101011101010100110101001101010001010011110100111101001111010100010101001101010101010101010101010101010101010101010101010101010101010101010101000110000111111101111110111110110111100000110111000111110111110111110111110,
	240'b101101001111111111101111101011101010011110101110110000111100111011001100110010001011111010110011101010111010011110101001101010101010101010101010101010101010101010101010101010001100101111111101111101001100111110111010111110111110111110111110,
	240'b101101001111111111101111101011001011101011101010111111011111111111111111111111111111110011110101111001011100111010110101101010011010100010101010101010101010101010101010101010101010100011010110111111111110010010111001111110111110111110111110,
	240'b101101001111111111101101101110101111000111111111111111111111111111111111111111111111111111111111111111111111111111110110110110101011011010101000101010011010101010101010101010101010100110111100110110101100100010111001111110111110111110111110,
	240'b101101001111111111101101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111001101101010111010100110101010101010101010101010101010101010011010011110111001111110111110111110111110,
	240'b101101001111111111110100111101101111111111111111111111111111111111111111111111111111111011111110111111101111111011111101111111111111111111111110110111111011000110101000101010101010101010101010101010101010100010111001111110111110111110111110,
	240'b101101001111111111111000111111001111111111111111111111111111111111111111111111001100111011000100110001011100010011100010111111111111111111111111111111111110101010110100101010001010101010101010101010101010100010111001111110111110111110111110,
	240'b101101001111111011111001111111001111111111111111111111111111111111111111111110101011010110100101101001101011001111110100111111111111111111111111111111111111111111101011101100111010100010101010101010101010100010111001111110111110111110111110,
	240'b101101001111111111110111111110111111111111111111111111111111111111111111111110101011011110101000101010101010110011011000111111111111111111111111111111111111111111111111111001101010111010101001101010101010100010111001111110111110111110111110,
	240'b101101001111111111110101111110011111111111111111111111111111111111111111111110101011011010100110101010101010100110101100110111101111111111111111111111111111111111111111111111111101100010101001101010101010100010111001111110111110111110111110,
	240'b101101001111111111110010111100101111111111111111111111111111111111111111111110011100001011000101101010101010101010101001101011111110010111111111111111111111111111111111111111111111110011000010101010001010100010111001111110111110111110111110,
	240'b101101001111111111101110111001111111111111111111111111111111111111111111111110111110110111110101110010101010100010101010101010001011001011101011111111111111111111111111111111111111111111101100101011101010011110111001111110111110111110111110,
	240'b101101001111111111101100110101101111111111111111111111111111111111111111111111111110101010111110111011001100010010100111101010101010100010110110111100011111111111111111111111111111111111111111110011001010011010111001111110111110111110111110,
	240'b101101001111111111101101110001001111110111111111111111111111111111111111111111111101001110100100101111111110110110111101101010001010101010100111110000011111101111111111111111111111111111111111111011101010110010111000111110111110111110111110,
	240'b101101001111111111101110101100111111000011111111111111111111111111111111111111111100110110100111101001111100010111101011101110001010100010101010101010111110101011111111111111111111111111111111111111101100001010110111111110111110111110111110,
	240'b101101001111111111101111101011001101011111111111111111111111111111111111111111111101011110100111101010101010100011001100111010011011001110101000101010011101111011111111111111111111111111111111111111111101110110111000111110111110111110111110,
	240'b101101001111111111101111101011001011101011111011111111111111111111111111111111111111000010110001101010001010101010101001110101001110010110101111101001111110001111111111111111111111111111111111111111111111000111000000111110101110111110111110,
	240'b101101001111111111101111101011101010100111100001111111111111111111111111111111111111111111011110101011001010100110101001101010101101101011011110101101101111010011111111111111111111111111111111111111111111110011001110111110011110111110111110,
	240'b101101001111111111101111101011101010011110111011111110101111111111111111111111111111111111111111110101111010101010101001101010011010110011011111111100101111001111111110111111111111111111111111111111111111111111011110111110011110111110111110,
	240'b101101001111111111101111101011101010100110101001110101111111111111111111111111111111111111111111111111101101000010101000101010101010100110110001110100001100110111111111111111111111111111111111111111111111111111101100111110011110111110111110,
	240'b101101001111111111101111101011101010100110101001101100001110110111111111111111111111111111111111111111111111110011001001101010001010101010101001101001101100010111111111111111111111111111111111111111111111111111110100111110111110111110111110,
	240'b101101001111111111101111101011101010100110101010101010001011101111110111111111111111111111111111111111111111111111111001110000111010100110101010101001111100011011111111111111111111111111111111111111111111111111110111111111001110111110111110,
	240'b101101001111111111101111101011101010100110101010101010101010100011000101111110101111111111111111111111111111111111111111111010011010101110100111101001011100010111111111111111111111111111111111111111111111111111111001111111011110111110111110,
	240'b101101001111111111101111101011101010100110101010101010101010101010101000110001111111100011111111111111111111111111111101110101001011101110111011101110011101001011111111111111111111111111111111111111111111111111111001111111011110111110111110,
	240'b101101001111111111101111101011101010100110101010101010101010101010101010101010001100000111110010111111111111111111111110111110101111101111111011111110111111110011111111111111111111111111111111111111111111111111110100111110111110111110111110,
	240'b101101001111111111101111101011101010011110101000101010101010101010101010101010101010100010110110111000001111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111110011110111110111110,
	240'b101101001111111111101110101100011100101111010000101101001010100110101010101010101010101010101000101010111100010011101001111111101111111111111111111111111111111111111111111111111111111111111111111111111110100110111111111110101110111110111110,
	240'b101101001111111111101110101101011111010011111110110000101010011110101010101010101010101010101010101010101010100010101101110000111110000011110010111111101111111111111111111111111111111111111111111010111011011010110111111110111110111110111110,
	240'b101101001111111111101110101101011110001011111101111100011011011110101000101010101010101010101010101010101010101010101001101010001010100110110010101111101100110011010110110110111101100111001000101011111010011010111001111110111110111110111110,
	240'b101101001111111111101111101100001100100011100001111111111110101110110010101010011010101010101010101010101010101010101010101010101010101010101001101010001010100010101000101001111010011110101000101010011010100010111001111110111110111110111110,
	240'b101101001111111111101110101011101110011111101001111000101111111111011001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111110111110111110111110,
	240'b101101001111111111101111101011011101100011111111111000111110100111100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111110111110111110111110,
	240'b101101001111111111101111101011011011000111101010111111111110000111000111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111110111110111110111110,
	240'b101101001111111111101111101011101010011110110110111011111111110111100100101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111110111110111110111110,
	240'b101011111111111111110011101100001010100110100111110000101111111111110011101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111100111111011110111110110110,
	240'b100111101111010011111110110010001010011010100110101100001100010111000000101010011010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010100011011000111111111110001110011011,
	240'b101110011101010111111111111101111101001111000101110001011100001111000100110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101101101011111100111111111100011010110111,
	240'b111011001011100111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100001011101100,
	240'b111110001110110010111100110101001110111111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110111110101011001110110001001111001111111000,
	240'b111111111111111111100101101000001001110010110001101100111011001110110011101100111011001110110011101100101011001010110010101100101011001110110011101100111011001110110011101100111011001010110011101011011001011110110110111110111111111111111111,
	240'b111100011111010011101100101010101010010110101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011011010001010101110111011001111001011110001,
	240'b111100001110101011000101110010011110001111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100001101110111000001110001011110111111110000,
	240'b111011111011110111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101100100011110000,
	240'b110000111100111011111111111101111011110110100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100001100111101001111010100001101000111100101011111110111111101100001011000011,
	240'b100111101111000111111110100111110101000101001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111101011000011110110111100101010111010011100101011110111110111111111101111110011011,
	240'b101011011111111111101011011000110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101111110011001100101010100100100111101111110111111001110111110110011,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110010111010011111111110111001010101100101000001110011111101101111000010111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000100110101101110011111111101010100101000101110010111101101111000010111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110110110001011110011100011111111011000010101101110111101101111000010111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111011111011110110101111011111010110101101101111101101111000010111110,
	240'b101101001111111111011111010111100101001101010011010100000100111101001111010100000101000101010011010101000101010101010101010101010101010101010101010101010101010101010010100001111111011111101110101101101000010001110000111101101111000010111110,
	240'b101101001111111111011111010111100101000001011110100010001001110110011010100100010111110001100110010101110101000001010010010101010101010101010101010101010101010101010101010100011001100011111011111010011001111101110101111101011111000010111110,
	240'b101101001111111111011111010110100111010111010101111111001111111111111111111111111111100011101100110010101001110101101011010100110101001001010101010101010101010101010101010101000101001010101101111111111100100101110011111101011111000010111110,
	240'b101101001111111111011100011101001110001111111111111111111111111111111111111111111111111111111111111111111111111111101100101101010110110101010001010101000101010101010101010101010101001001111001101101101001000101110011111101011111000010111110,
	240'b101101001111111111011100101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110011010010101110101001001010101010101010101010101010101010100100100111101110011111101101111000010111110,
	240'b101101001111111111101001111011101111111111111111111111111111111111111111111111111111110111111101111111011111110111111011111111111111111111111110101111110110001001010001010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111110001111110011111111111111111111111111111111111111111111110001001110010001000100010101000100111000100111111111111111111111111111111111101010001101001010100010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111110010111110011111111111111111111111111111111111111111111101010110101001001101010011010110011111101010111111111111111111111111111111111111111111010111011010000101000101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111101111111110001111111111111111111111111111111111111111111101010110111001010010010101000101100010110001111111111111111111111111111111111111111111111111110011010101110101010011010101010101000101110011111101101111000010111110,
	240'b101101001111111111101011111101001111111111111111111111111111111111111111111101010110110001001110010101010101001101011000101111011111111111111111111111111111111111111111111111111011000001010011010101000101000101110011111101101111000010111110,
	240'b101101001111111111100101111001011111111111111111111111111111111111111111111100111000010010001100010101000101010001010010010111111100101111111111111111111111111111111111111111111111100110000101010100000101000101110011111101101111000010111110,
	240'b101101001111111111011110110011111111111111111111111111111111111111111111111101111101101111101010100101010101000001010101010100010110010111011000111111111111111111111111111111111111111111011001010111010101000001110011111101101111000010111110,
	240'b101101001111111111011001101011101111111111111111111111111111111111111111111111111101010101111100110110011000100101010000010101010101000101101110111000101111111111111111111111111111111111111111100110010100110001110011111101101111000010111110,
	240'b101101001111111111011010100010001111101011111111111111111111111111111111111111111010011101001010011111111101101101111100010100000101010101010000100000111111100011111111111111111111111111111111110111000101101001110001111101101111000010111110,
	240'b101101001111111111011101011010001110000011111111111111111111111111111111111111111001101101001111010100001000101111010111011100010101000101010100010101111101010111111111111111111111111111111111111111011000011001101110111101101111000010111110,
	240'b101101001111111111011110010110101011000011111111111111111111111111111111111111111010111001001111010101000101000110011001110100110110011101010001010100101011111011111111111111111111111111111111111111111011101001110001111101011111000010111110,
	240'b101101001111111111011111010110100111010111110110111111111111111111111111111111111110000101100010010100100101010001010011101010001100101001011111010100001100011011111111111111111111111111111111111111111110010010000001111101001111000010111110,
	240'b101101001111111111011111010111010101001111000011111111111111111111111111111111111111111110111110010110010101001101010100010101101011011010111101011011011110100111111111111111111111111111111111111111111111100010011101111100011111000010111110,
	240'b101101001111111111011111010111100100111101111000111101011111111111111111111111111111111111111111101011110101010001010100010100110101101010111110111001001110011011111101111111111111111111111111111111111111111110111101111100011111000010111110,
	240'b101101001111111111011111010111100101001101010010101011111111111111111111111111111111111111111111111111011010000101010010010101000101001001100100101000011001101111111110111111111111111111111111111111111111111111011001111100101111000010111110,
	240'b101101001111111111011111010111100101001101010011011000011101101111111111111111111111111111111111111111111111100010010011010100010101010101010100010011011000110111111111111111111111111111111111111111111111111111101010111101001111000010111110,
	240'b101101001111111111011111010111100101001101010101010100010111100011101110111111111111111111111111111111111111111111110011100010000101001101010101010100001000111011111111111111111111111111111111111111111111111111101111111101111110111110111110,
	240'b101101001111111111011111010111100101001101010101010101010101000010001100111101001111111111111111111111111111111111111111110101000101100001001111010011001000101111111111111111111111111111111111111111111111111111110010111110011110111110111110,
	240'b101101001111111111011111010111100101001101010101010101010101010001010001100011111111001011111111111111111111111111111011101010010111011001111000011101001010011011111111111111111111111111111111111111111111111111110010111110011110111110111110,
	240'b101101001111111111011111010111100101001101010101010101010101010101010100010100011000001111100110111111111111111111111101111101011111011011110111111101101111100111111111111111111111111111111111111111111111111111101000111101001111000010111110,
	240'b101101001111111111011111010111100100111101010000010101000101010101010101010101010101000101101100110000011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010111100011111000010111110,
	240'b101101001111111111011110011001001001011010100010011010000101001101010101010101010101010101010001010101111000101011010011111111001111111111111111111111111111111111111111111111111111111111111111111111111101001101111110111101001111000010111110,
	240'b101101001111111111011101011010101110100111111110100001010100111101010101010101010101010101010101010101000101000001011100100001111100000111100110111111001111111111111111111111111111111111111111110101100110110101101111111101101111000010111110,
	240'b101101001111111111011101011010101100011011111011111001000110111001010001010101010101010101010101010101010101010101010100010100000101001101100101011111101001100010101100101101101011010010010000010111110100111001110011111101101111000010111110,
	240'b101101001111111111011110011000001001000011000010111111111101100001100110010100110101010101010101010101010101010101010101010101010101010101010011010100010101000001010000010100000101000001010000010100110101000101110011111101101111000010111110,
	240'b101101001111111111011110010111011100111111010100110001101111111110110011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111011110010110111011000111111111110001111101001011001000010101010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111011111010111000110001111010110111111111100010010001110010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101101001111111111011111010111100100111101101101110111111111110011001001010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101101111000010111110,
	240'b101011111111111111100111011000010101001101001111100001001111111111100110010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001111001111110101111000010110110,
	240'b100111101111010011111100100100010100111001001101011000011000110010000001010100100100111101010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110101000110110000111111111110001110011011,
	240'b101110011101010111111111111100001010011010001100100011001000100010001001100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011011011011111010111111111100011010110111,
	240'b111011001011100111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100001011101100,
	240'b111110001110110010111100110101001111000011111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110101011001110110001001111001111111000,
	240'b111111111111111111100101101000001001110010110001101100111011001110110011101100111011001110110011101100101011001010110010101100101011001110110011101100111011001110110011101100111011001010110011101011011001011110110110111110111111111111111111,
};
assign data = picture[addr];
endmodule