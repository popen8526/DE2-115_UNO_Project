module red_two(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
    240'b111101001111110011010111101101101011011110111000101110001011100010111000101110001011100010111001101110011011100110111001101110001011100010111000101110001011100010111000101110011011100110111001101110001011010110110100110101011111000111110000,
    240'b111101111101010011001000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111101101000111110011,
    240'b110101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011110011011110,
    240'b101100011111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010101011,
    240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010100110,
    240'b101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
    240'b101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010,
    240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010100100,
    240'b101101011110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010110011,
    240'b111000001100000111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011100111100110,
    240'b111101111101110111000001111011001111100111111001111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110011111100111100110101110011101101011110011,
    240'b111110001111011111011000100011101001010110101100101011001010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100101010101001000010011100111010011111111011111010,
    240'b111101001111110011010111101101101011011110111000101110001011100010111000101110001011100110111001101110011011100110111001101110001011100010111000101110001011100010111001101110011011100110111001101110001011010110110100110101101111001011110000,
    240'b111101111101010011001000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111101101000111110011,
    240'b110101111100011111111111111111111111001111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100110111001111111011111111111111110111011110011011110,
    240'b101100011111001011111111110001010111010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110001001100100011000100111101111010110111111111110011010101011,
    240'b101101011111111111100111011001010100111101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010010010101101001010110111100100101000101000101110101111101011111110110100110,
    240'b101110111111111111000110010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101001001111011111011011111101111010000101011000110111011111111110110011,
    240'b101111001111111111000001010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111000101010101001010011101011101110010001100011110101111111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111001101001110001001010011010011000101101100001110110001111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101100101110101101111111010011100100111001011011110110011111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010001010100010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010110001011100111110010101000010101011101011010110110011111111110110101,
    240'b101111001111111111000001010101000101001101010001010100110101100001010111010100110101000001010000010100100101010001010101010101010101010101010101010101010101010001011011100010110110111110101100111110101011101001100000110110001111111110110101,
    240'b101111001111111111000001010100100101010110000110101111101100111011001100110001011011000010010010011100010101100101010000010100110101010101010101010101010101001101100011111011011110010011010100111110111110110101101011110101111111111110110101,
    240'b101111001111111111000000010101101010111111111001111111111111111111111111111111111111111111111111111100011101000110011000011000100101000001010011010101010101010001011101101010001011100010111000101101101010010001100011110110001111111110110101,
    240'b101111001111111110111110100110011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111000001001011001011011010100010101010101010101010100100101001001010010010100100101000101011011110110011111111110110101,
    240'b101111001111111111001110111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001101011100110101000101010100010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111100100111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000100101010001010101000101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111101110111111001111111111111111111111111111111111111111111111111111111111111111111111111111011011011000110011001101110111111011111111111111010110010100010100010101010001010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111101101111111001111111111111111111111111111111111111111111111111111111111111111110100010111110001011000010100110101110010001001111000001111111111110110100011110101000101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111101001111110111111111111111111111111111111111111111111111111111111111111010001011000010100111001001111010011110100111101001110011011111110010011111111111100000111110001010001010101010101010001011011110110011111111110110101,
    240'b101111001111111111100010111110011111111111111111111111111111111111111111111111111111011001111010010011100101100110010010101011111000010101010101010011101001001111111101111111111101110101100100010100100101010001011011110110011111111110110101,
    240'b101111001111111111010111111011101111111111111111111111111111111111111111111111111101000001010110010100101010011111111110111111111111011110001110010011110110001111100111111111111111111110110100010100110101001101011011110110011111111110110101,
    240'b101111001111111111001001110110111111111111111111111111111111111111111111111111111011001101001110011000111110100011111111111111111111111111001111010100000100111111001110111111111111111111110111011111000100111101011011110110011111111110110101,
    240'b101111001111111110111110101111001111111111111111111111111111111111111111111111111010111101001101011001101110110111111111111111111111111111101000100100011000110011011010111111111111111111111111110010000101010101011010110110011111111110110101,
    240'b101111001111111110111100100100111111111111111111111111111111111111111111111111111100010101010011010101011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111100101010111110110011111111110110101,
    240'b101111001111111110111110011010101110111111111111111111111111111111111111111111111110110001101001010011100111000011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111011010101011000110110011111111110110101,
    240'b101111001111111111000001010100111100001111111111111111111111111111111111111111111111111110111011010101110100111101101010110010111111111111111111111111111111111111111111111111111111111111111111111111111110010001101000110101111111111110110101,
    240'b101111001111111111000001010011111000010111111100111111111111111111111111111111111111111111111110101101000101100101001111010111001010101111110110111111111111111111111111111111111111111111111111111111111111110010001011110101001111111110110101,
    240'b101111001111111111000001010100110101100111010000111111111111111111111111111111111111111111111111111111111011111101011111010011110101001010000011111000011111111111111111111111111111111111111111111111111111111110110001110101001111111110110101,
    240'b101111001111111111000001010101000101000010000011111110101111111111111111111111111111111111111111111111111111111111010010011100110101000001001111011010001100001111111100111111111111111111111111111111111111111111010001110110101111111110110101,
    240'b101111001111111111000001010101000101010001010100101110101111111111111111111111111100010110000101100110101111100111111111111011001001000101010110010100010101101011010011111111111111111111111111111111111111111111100111111000101111111110110101,
    240'b101111001111111111000001010101000101010001010010011001101110000111111111111111111010011101001000010110001001001010010111100110101001000001011110010100110101001111000110111111111111111111111111111111111111111111110101111010101111111110110101,
    240'b101111001111111111000001010101000101010001010101010100010111110111110001111111111010100101001101010100110100111101001111010011110101000001010011010100100101001011000110111111111111111111111111111111111111111111111001111011101111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101000110001110111110001011001101011001010111110101111101011111010111110101111101011111010111100101111011001010111111111111111111111111111111111111111111111010111100011111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010001100100101110001111011110110111001101110011011100110111001101110011011100110111001101110011110100111111111111111111111111111111111111111111111010111100001111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010100010100011000010111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111010001111111110110101,
    240'b101111001111111111000001010101000101001101010100010101000101010001010100010101010101000101101110110000111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001110110011111111110110101,
    240'b101111001111111111000001010101010101100001011001010110010101100101011000010101010101010101010010010101111000101111010101111111001111111111111111111111111111111111111111111111111111111111111111111111111110111101111101110101011111111110110101,
    240'b101111001111111110111111011010111100011011010000110100101101001110110001010101110101010001010101010101000101000001011100100001111100000011101000111110101111111111111111111111111111111111111111111001101000011001011000110110011111111110110101,
    240'b101111001111111110111110011101011111110111101110101111101101110111010100010110000101010001010101010101010101010101010100010100000101010001100100100000011001100110101110101110001011101010011110011010100101000001011011110110011111111110110101,
    240'b101111001111111111000000010110111011100011110101101010100110100101101111010101100101010101010101010101010101010101010101010101010101010001010011010100000101000001010010010100110101001101010001010100100101010001011011110110011111111110110101,
    240'b101111001111111111000001010100100101010110011010111100101011110001011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111000001010100110100111001001111011111111110110110101000010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111110111111011001101010011001100101010010011011001011010110010101110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111110111110011001111111000010100100011001001101000011000110010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101110111111111111001001010100101010100111110111111011011110111101111111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011100111000001111111110110010,
    240'b101101001111111111101101011011010101000110001000101000010111010001001111010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100110110000010111110001111101110100100,
    240'b101101011110110011111111110101111000011101110011011100110111010101111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011101111001000111100101111111111110000010110011,
    240'b111000001100000111111010111111111111111011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111111111111111111101001011100111100110,
    240'b111101111101110111000001111011001111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011100110101110011101101011110011,
    240'b111110001111011111011000100011101001010110101100101011001010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100101010101001000010011100111010011111111011111010,
    240'b111101001111110011010111101101101011011110111000101110001011100010111000101110001011100010111001101110011011100110111001101110001011100010111000101110001011100010111000101110011011100110111001101110001011010110110100110101011111000111110000,
    240'b111101111101010011001000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111101101000111110011,
    240'b110101111100011111111111111111111111001111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100110111001111111011111111111111110111011110011011110,
    240'b101100011111001011111111110001010111010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110001001100100011000100111101111010110111111111110011010101011,
    240'b101101011111111111100111011001010100111101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010010010101101001010110111100100101000101000101110101111101011111110110100110,
    240'b101110111111111111000110010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101001001111011111011011111101111010000101011000110111011111111110110011,
    240'b101111001111111111000001010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111000101010101001010011101011101110010001100011110101111111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111001101001110001001010011010011000101101100001110110001111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101100101110101101111111010011100100111001011011110110011111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010001010100010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010110001011100111110010101000010101011101011010110110011111111110110101,
    240'b101111001111111111000001010101000101001101010001010100110101100001010111010100110101000001010000010100100101010001010101010101010101010101010101010101010101010001011011100010110110111110101100111110101011101001100000110110001111111110110101,
    240'b101111001111111111000001010100100101010110000110101111101100111011001100110001011011000010010010011100010101100101010000010100110101010101010101010101010101001101100011111011011110010011010100111110111110110101101011110101111111111110110101,
    240'b101111001111111111000000010101101010111111111001111111111111111111111111111111111111111111111111111100011101000110011000011000100101000001010011010101010101010001011101101010001011100010111000101101101010010001100011110110001111111110110101,
    240'b101111001111111110111110100110011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111000001001011001011011010100010101010101010101010100100101001001010010010100100101000101011011110110011111111110110101,
    240'b101111001111111111001110111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001101011100110101000101010100010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111100100111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000100101010001010101000101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111101110111111001111111111111111111111111111111111111111111111111111111111111111111111111111011011011000110011001101110111111011111111111111010110010100010100010101010001010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111101101111111001111111111111111111111111111111111111111111111111111111111111111110100010111110001011000010100110101110010001001111000001111111111110110100011110101000101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111101001111110111111111111111111111111111111111111111111111111111111111111010001011000010100111001001111010011110100111101001110011011111110010011111111111100000111110001010001010101010101010001011011110110011111111110110101,
    240'b101111001111111111100010111110011111111111111111111111111111111111111111111111111111011001111010010011100101100110010010101011111000010101010101010011101001001111111101111111111101110101100100010100100101010001011011110110011111111110110101,
    240'b101111001111111111010111111011101111111111111111111111111111111111111111111111111101000001010110010100101010011111111110111111111111011110001110010011110110001111100111111111111111111110110100010100110101001101011011110110011111111110110101,
    240'b101111001111111111001001110110111111111111111111111111111111111111111111111111111011001101001110011000111110100011111111111111111111111111001111010100000100111111001110111111111111111111110111011111000100111101011011110110011111111110110101,
    240'b101111001111111110111110101111001111111111111111111111111111111111111111111111111010111101001101011001101110110111111111111111111111111111101000100100011000110011011010111111111111111111111111110010000101010101011010110110011111111110110101,
    240'b101111001111111110111100100100111111111111111111111111111111111111111111111111111100010101010011010101011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111100101010111110110011111111110110101,
    240'b101111001111111110111110011010101110111111111111111111111111111111111111111111111110110001101001010011100111000011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111011010101011000110110011111111110110101,
    240'b101111001111111111000001010100111100001111111111111111111111111111111111111111111111111110111011010101110100111101101010110010111111111111111111111111111111111111111111111111111111111111111111111111111110010001101000110101111111111110110101,
    240'b101111001111111111000001010011111000010111111100111111111111111111111111111111111111111111111110101101000101100101001111010111001010101111110110111111111111111111111111111111111111111111111111111111111111110010001011110101001111111110110101,
    240'b101111001111111111000001010100110101100111010000111111111111111111111111111111111111111111111111111111111011111101011111010011110101001010000011111000011111111111111111111111111111111111111111111111111111111110110001110101001111111110110101,
    240'b101111001111111111000001010101000101000010000011111110101111111111111111111111111111111111111111111111111111111111010010011100110101000001001111011010001100001111111100111111111111111111111111111111111111111111010001110110101111111110110101,
    240'b101111001111111111000001010101000101010001010100101110101111111111111111111111111100010110000101100110101111100111111111111011001001000101010110010100010101101011010011111111111111111111111111111111111111111111100111111000101111111110110101,
    240'b101111001111111111000001010101000101010001010010011001101110000111111111111111111010011101001000010110001001001010010111100110101001000001011110010100110101001111000110111111111111111111111111111111111111111111110101111010101111111110110101,
    240'b101111001111111111000001010101000101010001010101010100010111110111110001111111111010100101001101010100110100111101001111010011110101000001010011010100100101001011000110111111111111111111111111111111111111111111111001111011101111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101000110001110111110001011001101011001010111110101111101011111010111110101111101011111010111100101111011001010111111111111111111111111111111111111111111111010111100011111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010001100100101110001111011110110111001101110011011100110111001101110011011100110111001101110011110100111111111111111111111111111111111111111111111010111100001111111110110101,
    240'b101111001111111111000001010101000101010001010101010101010101010101010100010100011000010111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111010001111111110110101,
    240'b101111001111111111000001010101000101001101010100010101000101010001010100010101010101000101101110110000111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001110110011111111110110101,
    240'b101111001111111111000001010101010101100001011001010110010101100101011000010101010101010101010010010101111000101111010101111111001111111111111111111111111111111111111111111111111111111111111111111111111110111101111101110101011111111110110101,
    240'b101111001111111110111111011010111100011011010000110100101101001110110001010101110101010001010101010101000101000001011100100001111100000011101000111110101111111111111111111111111111111111111111111001101000011001011000110110011111111110110101,
    240'b101111001111111110111110011101011111110111101110101111101101110111010100010110000101010001010101010101010101010101010100010100000101010001100100100000011001100110101110101110001011101010011110011010100101000001011011110110011111111110110101,
    240'b101111001111111111000000010110111011100011110101101010100110100101101111010101100101010101010101010101010101010101010101010101010101010001010011010100000101000001010010010100110101001101010001010100100101010001011011110110011111111110110101,
    240'b101111001111111111000001010100100101010110011010111100101011110001011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111111000001010100110100111001001111011111111110110110101000010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111110111111011001101010011001100101010010011011001011010110010101110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101111001111111110111110011001111111000010100100011001001101000011000110010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110011111111110110101,
    240'b101110111111111111001001010100101010100111110111111011011110111101111111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011100111000001111111110110010,
    240'b101101001111111111101101011011010101000110001000101000010111010001001111010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100110110000010111110001111101110100100,
    240'b101101011110110011111111110101111000011101110011011100110111010101111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011101111001000111100101111111111110000010110011,
    240'b111000001100000111111010111111111111111011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111111111111111111101001011100111100110,
    240'b111101111101110111000001111011001111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011100110101110011101101011110011,
    240'b111110001111011111011000100011101001010110101100101011001010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100101010101001000010011100111010011111111011111010,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule