module Background(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 600;
localparam Y_WIDTH = 430;
localparam [0:85][959:0] r_picture = {
	960'b000010110000101100001100000011100000111100001111000011100001000100010011000100110001001000010001000100100001000100010010000100010001001000010100000100110001001000010000000100000001000100010000000100010001000000010001000100110001001100010010000100000001000100010001000100000001000100010000000100100001001100010011000100100001000000010001000100000001000100010000000100000001001000010010000100100001000000001110000100000001000000010001000011110001000000010010000100100001000100010000000011110001000000001111000100000000111100010010000101000001010000010010000100000001000000001111000011110000111100001111000100010001001000010010000100010001001000010010000100000001001000010000000100000001010000010011000100100001001000010010000100010001000100010010000100100001001100010100000100110001000100010001000100100001000000010001000100010001000000010010000101000001001100001111000100000001001000010000000100100001000100010000000100100001000100010000000011010000110100001110,
	960'b000010110000110100001110000011110001000100010100000101000001010100011000000101100001010100011000000101010001001100010101000101110001010000010111000110000001010000010100000101100001010000010011000101010001010100010010000101110001011000010011000101010001011100010100000101000001010100010100000100110001011100010111000101000001010100010110000101000001010100010110000100110001010100011000000101010001001100010110000101010001001100010101000101100001001100010101000101010001010000010100000101110001010000010010000101010001010100010011000101100001011100010100000101000001011000010010000100100001011000011000000101100001011100010110000101000001011000010100000101000001010100010111000101000001011000010110000101010001011100010110000101000001010000010110000101100001010000011000000101100001001100010110000101010001010000010100000101010001010000010011000101100001010100010011000101010001010000010011000101000001011000010101000101000001010100010100000100100000111100001110,
	960'b000011000000111000010000000101000001010100010110000110100001100000011011000110010001110000011001000110100001110100011010000110110001110000011000000110110001100100011101000110010001101100011101000110010001101000011011000110000001100100011000000111000001100000011011000110110001100100011100000110010001100100011001000110100001100100011001000110110001101000011001000110100001100000011011000101110001101100011001000101110001110000011000000110000001101100010111000110010001011100011011000110100001100000011000000110010001100100011010000110010001100100011000000110110001100000011001000110000001011100011001000110000001101000011000000110000001100100011011000111010001100000011010000111000001100100011001000110110001101100011000000111010001110100011000000110110001101000011010000110010001101100011010000110010001110000011010000110100001110000011001000110100001011100011011000110010001100100011100000110100001101000011011000110000001100000010110000101100001001000010000,
	960'b000011100000111100010010000101110001100000011001000111000001111000011100000111110010000000011110000111110010000100011101000111100001111100011110000110110001111000011110000111000001111100100010000111110001111100100010000111110001110100100000000111010001110000100000001000000001110000011101001000010001110000011101001000000001110100011101001000010001111100011110000111100001111000011011000111100001111100011101000111100010000100011101000110100010000000011110000110100001110100011101000110110001110100100000000111010001110000100000000111010001110100011111000111000001110100011110000111110001110000011100000111100001101100011011000111000001111000011111001000000001111000011100000111100001110000011101000111110001110100100000001000000010000000011110000111100001111100011100000110110001111000011100000111100010000100011110000111100001111100100000000111000001111000011110000111010001110100100001000111100001110000011111000111010001101000011011000110000001011000010011,
	960'b000011100001010000011001000110010001110100100001000111110001111100100010001000000010000000100100001000110010000100100101001001010010000000100000001000100001111100011111001001000010001100100011001001010010001100100000001000010010000000100000001000010010010100100011001000100010010000100000000111110010001000100000000111110010001000100100001000100010010000100100001000010001111100100000000111110001111100100100001000110010001100100100001000100010000000011111001000010001111100100001001001000010001000100000001000110010001100011111001000000010000100100000001000100010010000100010001000110010011000100010000111110010000000011111000111000010001000100100001000100010011000100010001000000010000000100010000111100010000100100101001000110010010000100110001000100001111100100001001000010001111100100011001001010010001000100100001001010010000000100000001000110001111100011111001001000010010000100000001001010010001100011110000111100010000000011100000110010001101100010110,
	960'b000100010001010000011001000111010001110100100000001000010010001100100001001001000010010000100100001000100010011000100101001001010010010000100001001000010010010000100100001001100010001100100101001001010010010000100101001000110010001100100100001000100010010100100100001001000010001100100011001001010010001000100011001000110010001000100010001001010010010000100100001000110010001100100001001000100010010000100101001001010010011000100101001000100010001000100011001000110010010100100101001001010010010000100110001000110010001100100110001000110010001100100110001001010010001100100101001001010010011000100011001001000010001000100010001000110010001000100110001001100010001100100011001001100010001000100011001001000010001100100011001001100010010100100100001001000010010100100010001001000010011000100100001001000010011000100011001000110010001100100100001000110010001100100101001000100010001100100111001001000010001000100011001000100001111100100010000111010001101000011000,
	960'b000101000001010100011001001000110010000000011111001001000010010000100101001001010010100100100100001001100010101100100110001001110010100000100101001001100010010000101000001001010010011000101001001000110010011100101001001001100010011000100110001001110010010100101000001010000010001000101000001010000010011000100101001010010010010100100011001010100010100000100101001001110010001100100100001001000010011100100011001001010010100100100101001001000010011000100100001001000010001000100111001000110010011100101010001001010010010100100111001001000010010100100110001001100010001100101001001010000010010000100110001001100010010100100101001001100010010000100110001010000010001100101000001001010010001100100110001001100010100000100100001010000010011100100101001010010010010100100110001001010010101000100111001001010010100000100101001000110010100100100100001001010010010100101001001010000010011000101010001001010010001100100111001000110010001100100010001000100001101000011010,
	960'b000100110001100000011010001000000010000100100101001001010010010100101010001001110010100000101010001001110010100000100110001010110010100000101001001010100010100000101010001010100010011000100111001001110010101100101001001010010010100100100110001010010010100000100111001010000010100000101010001001110010101000101000001010100010101100100110001001110010010100101010001010100010011100101010001010000010100000101000001001010010011100100111001010110010100000101001001010100010001000100111001010000010010100100110001001100010100000100111001001110010100100100101001001110010011100100101001001010010100000100111001001010010100100101001001001110010101000100101001001100010100100101010001001010010101100101101001001010010100100101010001001110010011100101010001010000010011100101101001010110010100000101010001010010010010100100110001010100010100000101001001011000010101000100111001011000010100000100110001010000010101000101000001010010010100100100011001000010001111100011010,
	960'b000100100001011100011101000111100010001100100100001001010010100100101100001011010010011000101010001010100010011100101011001010010010100000101010001010010010101000101001001010000010101100100111001010110010100000101000001011100010110000101000001001110010101000101010001010010010101100101000001010010010110100101100001010010010101000101100001001110010100100101010001010000010101100101100001010110010100000101001001010100010011100101011001010000010011000101101001011000010100100100110001010100010101100100111001010010010011000100110001011000010110100101001001001110010101000101000001010000010101000100110001010000010110000101100001001110010101000101000001010000010100100100111001010010010110000101100001010100010011000101010001001110010100000101001001010000010100100101010001010100010101000100111001010010010100000101011001010010010100000101010001011000010101100101001001010000010101000100111001010100010100000101000001010010010100100100110001000000001111000011011,
	960'b000101100001011100011011001000000010001000100101001010100010101100101101001011000010111100101010001001110010100100101000001011010010111100101011001010010010110100101110001010100010100100101010001010010010100100101111001011010010101100101110001011100010100100101010001010010010100100101101001011100010101100101011001011110010101000101010001010000010100100101001001011100010101100101010001010100010111100101001001001110010100100101000001010000010111000101010001010110010110000101111001010100010100100101001001001110010100100101110001010010010100100101011001010110010011100100111001001110010100100101100001010110010101100101010001011000010101000101000001010100010100100101110001011110010110000101101001011110010110100100111001010000010100100101011001100010010111000101101001011000010111000101101001001110010101100101000001010100010111100101110001011000010110100101111001011000010101000101100001010000010110000101111001010100010100000100110001001000001111100011001,
	960'b000101010001011000011100000111110010001000100101001010010010101000101100001010110010110000101000001001110010100100101001001010100010110100101100001010100010101100101011001010000010100100101001001010000010101000101100001010100010101100101110001011010010100000101010001010010010100000101100001011000010101000101011001011010010101000101001001010100010100100101000001011010010101100101011001010100010110100101000001010010010101000101001001010010010111000101010001010110010100100101101001010000010100000101000001010000010100100101100001010110010100100101001001010000010100100101001001010010010100000101010001010100010101100101001001010110010101000101001001010010010101000101000001011100010110000101101001011000010101000101001001010000010100100101000001011000010101100101100001010110010110000101000001010100010101000101001001010100010101100101100001011000010110000101110001010010010100100101001001010100010011100101110001010100010100000100111001000110001111000011011,
	960'b000100100001100100011110000111100010001100101000001001100010110000101110001011100010100100101100001011000010011100101010001010110010011100101111001011100010110100101001001011000010100100101001001011000010100100101010001011010010110100101001001001100010101100101000001010000010101000101000001010000010110000101010001001110010100100101010001001110010100100101001001010000010101100101101001011010010011100101010001010110010011000101010001010000010100000101110001011000010101000100110001010010010011100100110001010110010100100101001001011010010110000101000001010000010100100100111001001100010100000101000001010100010111100101110001001110010110100101011001010000010101100101011001010010010110100101101001010010010100000101010001010000010100100101010001010010010101100110000001011100010100100101100001011010010100000101011001011100010100100101100001011110010111100100110001010110010101100100110001010110010101100100111001011010010110100100101001000100010001000011101,
	960'b000101000001101000011101001000000010001000101000001010010010100100101110001010100010100100101001001010100010111000101000001010110010101100100111001011010010100000101101001011010010100100100110001000100010010100100101001010010010101100101011001011000010110000101010001010100010110000101011001010100010110100101010001010100010101100101010001010110010100100101011001011000010101000101110001010000010011100101010001001100010011100100101001001110010010100100111001010000010011000100111001001110010011000100101001001100010100000100101001001100010100000100111001010000010011100101000001011000010101100101011001010110010110000101010001010010010101100101011001010110010101100101100001010110010101000101010001010100010100100101001001011010010101100101000001010000010001100100101001000110010100100101101001010010010110100101010001010110010111000101011001011100010100000101011001010110010100100101010001010010010101100101100001001110010100100100110001001000001111100011110,
	960'b000101100001011100011100001001010010001000100011001010100010101000101001001010110010101000100101001011010011001000101010001010100010110000101011001011000010101000100111001000000010101000111101010100100110000001100110011010100111000001110010011100010110111001101101011010110110010101100001010111100101111001011011010101100101010001010011010100100101010001010010010101000101010101010010100010101000111110010000100101101001111010100001101010101010111110110011101101101011011010110111101101101011011110110111101100111010111010101010101001001001111110010111100100001000110110000011010011110100110101001110010011110101000001010101010100110101001101010110010110010101101001011000010110110101111001100101011010010110110101101111011101010111101101110011011010110110011001011101010010110011010100100100001000100010100100101110001010110010110000101011001010010010101000101110001010110010101100110001001010110010100100101100001010000010011000100110001000110010000000011111,
	960'b000100110001100100011111001000110010001100101000001010000010101100100110001010010010100100101100001011100010111000101101001010110010101000101011001000100010010000111101011010101000001010000101011110110111001101110011011101100111011101110110011110100111111001111101011110100111011101110111011100110111001001110000011011000110100001100001010111100101110101011100010111100110000001011110011100001010111010110110101111011100100111010010110111001110011011101110111101011111100011111000111101111111011111110011111011011110011011011100110101001100101111000000101110011010100101101101010111110110000101100001011000110110010001100111011001010110011001101001011010100110110001101110011100010111010001111010011110110111110101111111100001001000100010000111100000111000001110000011100001011000011101111110010110100011001000100011001010100010100100101010001010010010100000101000001011000010111000101100001011000010110000101010001001100010011100100101001000110010001000011111,
	960'b000100010001100100100001001000000010010100101010001001010010011000101010001010100010100100101101001011100010111000101110001011000010010000100101010011000111110110001001100000100111000101110100011110010111111110000010011111110111111101111110011111010111110101111110011110110111011101110100011100110111000101110000011011110110101001100101011000010110001101100000011001000110010101100101010110110101111110000001100110001001111110100011101001101010100110101100101011101010111110110000101100001011000010101101101011001010100110100110101001001010000010011001100000010101111101100000011000100110001101100101011001010110001101100011011000010110010001100100011001010110100101101101011100000111011001111110100001001000100010001011100011101000110110001110100100101001010010010010100011011000011010000011100001111000010101101011001110100010001000100110001010110010101000101001001011010010110100101100001011100010110000101001001010000010011100100100001000100010001100011101,
	960'b000101010001011100011101001001010010000100100010001010000010100100101000001010110010110100101001001011000011000000101001001000100011111101111100100001010111010001110000011110011000000110000110100001111000011110000011100000111000000010000011100000101000001110000001100000101000000101111110011111000111101101110110011101010111000101110000011011110111001001110001011101000111001001110001011100010111010101101011011001010110011101100111011010000110100101100110011001010110010001100011011000110110010001100100011001000110010101100110011010000110011101101001011011010111001001110010011011110110111101110000011011110110111101101111011100000111010001110111011101110111100101111011011111101000000101111111100000111000001110000111100011111001001010010100100110001001011110011010100110011001010110001111100001010111101001111100100000000110010100110001001001010010101100101101001010100010101000101111001010100010011100101100001010000010010100100110001001010001111100011101,
	960'b000101000001100100011100001000100010001000100101001010110010100000101010001010100010110100101100001011010010100100101001011000101000000101110100011011100111011001111100100001111000110110010010100111101010111010111011110001111100110111001110110011111100111111001111110011111100111111001111110011111101000011010000110100001101000111010001110100011101001111010100110101001101010111010101110101011101010011010011110101001101010011010100110100111101010011010100110101001101010011010011110100111101001111010010110100101101001111010100110101001101010011010110110101101101010011010100110101011101010011010011110100011101000111010001110011111100111011001110110011001100110011001101110011111101000111010010110101001101010111010111110101111101011011010011110011001100000110110101101010001001111010010111100011011000011010000000011100010111011001111101010010000010001100101011001011010010101100101011001010010010110000101100001001100010100000100101001001010010000100011101,
	960'b000100100001100100011110000111110010010000101001001001110010101100110001001011000010100100101110001001010011001101110100011111010111001001111001011111101000010010001011101000011011111111010111111010001110111111101101111010001110001111100000111000001110000011100000111000001101111111011110110111011101111111011111110111111101111111100000111000011110000111100010111000111110001011100010111000111110001111100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001011110010011100100111001001110010011100101111001011110010111100101111001001110001111100011111000111110001011100001111000101110001011100001111000011110000111100010111000101110001011100010111000111110010011100100111001001110011011101000111011011111000011101111111001011101001110111000101000011001010010001100011111110111010101110010011111100110000100100111001001110010110000101000001011010010110100101000001011010010111000100101001000100010000100011110,
	960'b000101000001010100011101001000000010010000100101001010100010101100101100001011010010110000100010001111100111111110000001100000111000011110001011100011111010001111001100111010011111000011100100110100001011101010100111100111011001100110010111100101111001011110010110100101101001011010010110100101101001011010010111100101111001011010010110100110001001100010010111100101111001011110010111100101111001011010010110100101101001011110010111100101111001011110010111100101111001011010010110100101111001011110010111100101111001011010010110100101101001011010010101100101011001011010010110100101101001011010010111100101111001011110010111100101111001100010010111100101111001011110010111100101101001010110010111100101111001011110010111100101011001011010011001100111111010101110111110110101001110100011101101110111111011110110100000100100011000100110000011011110111000001101101100001010110010011000101001001010110010100100101110001010100010100100100111001001000001111000011100,
	960'b000101010001101000011101001000110010001000101000001011010010101100101100001010100010010101000100100001001000111110010011100110001010010110100101110001011110100011101111110101111011010110011010100001110111001001011111010011000100000100111101001110100011101000111100001111000011101100111011001110110011101000111011001110100011101000111010001110110011101100111011001110110011101100111011001110110011101100111010001110100011101000111010001110110011110000111100001111000011101100111101001111000011110100111101001111000011110000111011001111000011110000111100001110110011101100111010001110100011101000111011001110110011101100111011001110110011101100111011001110110011101000111011001110110011110000111100001111000011101100111011001110110011110001000100010100000110001001111000100011001001110110111011110111011110101111011001101100101001101010011111100101111000101010001000011100110010110100101000001010100010111000101111001010100010101000101000001001010010000000011101,
	960'b000100110001011100011111001000010010010100100100001010010010110000101111001001110011111110001100100111011010010010101111101110001011000111011000111011111101111110110000100011110110111101000010001000000000110000000101000001000000000100000011000000000000000100000001000000010000000100000000000000010000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000010000000000000001000000010000001000000010000000010000000100000100000000000000000000000000000000000000001000000001000000010000000000000001000000000000000100000000000000010000000100000000000000000000000100000001000000000000000000000000000000000000000000000001000000000000000000000000000000100000001000000010000000100000001100000010000000110000010100001111001001010100110001110100100100101011100011100001111001011100011010100010101010111010100110100000100101010111001100101010001010010010100000101010001011100010101100100111001000010001111100011111,
	960'b000100100001101000011110001000100010011000101010001010000010101000101000001101111000101010100001101100011100010011000011101111001110000111101011110000111001001001101001001100000000101000000010000000100000010000000100000001000000010000000100000000100000001100000010000000110000010000000011000000100000001000000010000000010000001000000001000000010000000100000010000000100000000100000001000000100000001000000010000000100000001000000010000000110000001100000011000000110000001100000011000001000000001100000010000000100000001100000011000000100000001000000010000000010000001000000001000000100000000100000001000000010000000100000010000000100000001000000000000000010000000100000001000000100000000100000010000000110000001100000001000000100000001100000011000000110000001100000100000000110000001000001111001110000110111110011011110010111110011011001110101001101011011010111001101010001001110001101000001001100010101000101011001010100010101100100100001001000010000100011100,
	960'b000101010001100000011101001001100010010100100100001010110010100000101010011111011010010010110010110011101100100110111101111001011110011110101111011110110011011100001001000000010000001100000011000000100000001000000011000000110000001100000100000000110000010000000011000000110000001100000011000000110000001100000100000000110000001100000011000000110000001100000011000000110000001100000100000000110000010000000100000000110000001000000011000000110000001100000011000000110000010000000100000000110000001100000100000000110000010000000011000001000000010000000100000000110000010000000011000000110000001000000011000000110000001100000100000000110000010000000011000000110000001100000011000000110000001100000011000001000000001100000011000000110000001100000100000000110000001000000100000000100000010000000100000000010000111001000101100000111011100111100010110011101010101011000001101110011010011110010100010101100010001100101100001001110010010100100101001001000001111000011110,
	960'b000101000001011100011101001000110010001000100011001010100010011001100000100111101010111011001010110011001011101111100110111000111010010001100001000110010000000100000100000000110000001100000011000001010000011000000101000001000000010000000011000000110000010000000011000000110000001100000011000001000000001100000011000001000000010000000100000001000000010000000011000001000000010000000011000001000000001100000011000001000000001100000011000001000000010000000100000001000000010000000100000000110000010000000100000000110000001100000100000001010000010000000011000001000000001100000011000000110000001100000100000000110000001100000100000000110000010000000100000001000000010000000100000001000000010000000011000001000000001100000011000000110000001000000100000001010000011000000101000001000000001000000011000001000000001100000011001001000110111110110000111000001100101010101001110001011011011110100011100001100011110100100111001010100010011100100111001000010010000000011111,
	960'b000100010001101000100001001000000010011100101010001000010100000010001001101001001011110011001101101100111110000011100101101000010101000100001011000000100000011000000011000000110000010100000101000000110000001000000010000000010000000100000001000000010000001000000001000000010000000100000001000000100000000100000010000000010000000100000010000000100000001000000010000000100000000100000010000000010000000100000001000000100000001000000010000000100000001000000001000000010000001000000010000000100000000100000001000000010000000100000010000000100000001000000001000000010000000100000001000000010000000100000010000000100000001000000010000000010000001000000001000000010000001000000011000000010000000100000001000000010000000100000010000000100000000100000010000000100000001000000010000001010000011100000100000000100000001100000101000000100001000101100001101011101101110111000000101010011100000110100111100011100110110000101010001001100010100000100011001000110010010000011111,
	960'b000100100001100000011110001000100010010000100100001001100110111010001001101000101100010110110001110101111110011110101000010010110000100100000100000001000000001100000100000001100000010000000010000000010000001000000010000000100000000100000001000000100000001000000010000000100000000100000001000000100000000100000001000000000000000100000001000000010000001000000010000000100000000100000001000000010000000100000001000000010000000100000010000000010000000100000010000000100000001000000010000000100000001000000001000000010000001000000010000000010000000100000001000000010000000000000001000000010000000100000011000000100000001000000010000000010000000100000001000000010000001000000011000000100000001000000010000000100000001000000010000000100000001000000001000000010000000100000001000000010000001000000110000001110000001100000011000000110000001000001100010111011011011011011001101101011010100010101110100100010111011101001011001001000010011100101000001000110010000000011101,
	960'b000101000001011100011100001001010010010100100001010011010111101110000111101010001010101111001001111001111011101001010010000010000000010000000101000000110000011000000101000000110000001100000001000000100000001000000010000000100000001000000010000000100000001000000010000000010000000100000001000000010000000100000010000000100000001000000010000000100000001000000010000000100000000100000001000000010000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000001000000010000000100000000100000000000000010000000100000001000000010000000100000001000000010000001000000010000000010000000100000001000000010000001100000011000000100000000100000010000000100000000100000001000000010000000100000010000000010000000100000010000000100000001000000010000000100000001000000010000000110000010100000100000000100000001100000010000011100110001111000100110011111010010110011111100100000111100001100000001100010010010100100110001000110001111000011101,
	960'b000100110001101000011100001000100010000100101100011010000111010110000100100110101011010011100100110100100110011100001110000001100000001000000011000001100000010000000010000000100000001000000010000000100000001000000001000000010000000100000010000000010000000100000010000000010000000100000001000000010000000100000001000000100000000100000001000000010000000100000001000000010000001000000010000000010000000100000001000000100000000100000010000000100000000100000010000000100000000100000001000000010000001000000011000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000100000001000000010000000010000000100000001000000010000000100000010000000010000000100000001000000100000001000000010000000100000000100000010000000010000000100000010000000110000001000000110000001000000001000000010000000100001010101111011110100101011111010010101100010100111011001100000010010010010011000100011001000110010001000011011,
	960'b000100110001011100011110001000010010000001001000011010100111000001111100100100011101001111100100100011100001110000000100000000100000001100000110000001000000000100000001000000010000000000000001000000010000000100000001000000100000000100000001000000010000000100000001000000010000000000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000110000001000000001000000100000000100000001000000010000000100000010000000100000000100000001000000010000000100000001000000000000000100000001000000010000000000000000000000010000000100000001000000010000000100000001000000010000000100000001000000100000000100000001000000110000001000000001000000100000000100000001000000100000001000000001000000000000000100000010000000010000001000000010000001100000010000000010000000110000001000101010101000101100111110100111100001010111010001100000010100010011000000100100001000000001110100011101,
	960'b000101110001100000011011001000000010011001011010011001010110100101110111101100011110000110111111001110100000001100000011000000100000010100000101000000110000001100000001000000100000000100000001000000010000001000000010000000010000000100000010000000100000000100000000000000010000000100000001000000010000000100000001000000100000000100000001000000100000001000000010000000010000000100000001000000010000000000000001000000010000001000000001000000100000001000000010000000100000000100000001000000100000000100000010000000100000001000000000000000010000000100000001000000000000000100000001000000000000000000000001000000010000000100000001000000100000000100000001000000100000001000000010000000100000001000000010000000100000000100000001000000100000000100000001000000100000001000000001000000010000001000000011000000100000001000000010000000100000011100000011000000110000010000000100010100011100011110111100100011110111001001100100010100010011111100100100001001010001111000011100,
	960'b000101100001100000011011000111010011100001011101011000010110001110000011110011001101111101110110000010110000010100000011000000110000011100000010000000110000001000000010000000110000001000000011000000100000001000000010000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000000000000100000010000000100000001000000010000000010000000100000010000000010000000100000001000000010000001000000001000000100000001000000010000000100000001000000001000000100000001000000010000000100000000100000001000000010000000100000001000000000000000100000001000000010000000100000001000000010000000100000001000000010000001000000010000000100000001000000010000000110000001000000010000000100000000100000001000000010000001000000001000000010000000100000010000000010000001000000011000000100000000100000001000000100000001100000110000000100000010000000011000100101001001111001001101000100111001101011111010100000100100100101000001000010001111000011101,
	960'b000100010001011100011110001000000100101101011000010110110110000010011111110110011100000000101101000000110000010100000100000001100000001000000001000000010000001100000011000000010000001000000011000000010000001000000001000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000100000000100000010000000100000000100000001000000010000001000000001000000010000000100000010000000010000000100000010000000010000000100000001000000010000000000000001000000010000000000000001000000010000001000000011000000010000000100000010000000100000000100000010000000010000000100000010000000100000001000000010000000010000000100000010000000100000000100000001000000010000001000000010000000100000001000000001000000010000000100000101000000110000001100000100000000110100011111000010101101001000000001011101010101010100011100110010001000000010000100011101,
	960'b000100100001100000011101001001010101010001010110010101100110110110110111110111001000011000001010000001000000010000000011000001010000000100000010000000100000001000000011000000100000000100000010000000010000001000000001000000010000000100000001000000010000000100000001000000010000001000000011000000100000001000000010000000100000000100000001000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000000000001000000010000000100000010000000000000000100000001000000010000000000000000000000000000000100000001000000110000000100000010000000010000000100000001000000100000000100000001000000010000000100000010000000100000001000000010000000010000000100000001000000100000001000000001000000100000001000000001000000010000001000000001000000010000001000000010000001100000001000000011000001000001010110011100101111111001001101100010010100110100010000111100001000000001111100011100,
	960'b000101010001011000011100001100100101010001010011010101100111111111000100110011110100010100000011000001000000001000000110000000110000001000000001000000110000001100000010000000100000000100000010000000010000000100000001000000010000000100000001000000100000001000000001000000010000001000000011000000100000000100000001000000100000000100000001000000100000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000000000000010000000100000001000000010000000100000010000000100000000100000001000000010000001000000001000000100000000100000001000000010000000100000001000000100000000100000001000000010000001000000001000000010000001000000010000000010000000100000010000000100000000100000010000000010000001000000010000001010000001100000010000001000000001101011110110000101010001001101011010101000100101001000001001001010001111000011110,
	960'b000100110001100000011101001111000100111101010001010110101001000111001000101011110001011100000100000001000000001000000110000000100000001000000010000000010000001100000010000000010000000100000001000000100000000100000001000000100000000100000001000000100000001000000010000000100000001000000010000000100000000100000010000000110000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000001000000010000000010000000100000000000000000000000100000001000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000001000000010000000010000000100000001000000100000000100000001000000100000000100000001000000010000000100000010000000100000000100000010000000010000000100000011000000110000010100000100000000110000001100101011101101111010110101110111010101010100110101000010001010000010000100011110,
	960'b000100100001101100100001010000010100110001010010011000011001110111001010100000110000010100000101000000110000010000000101000000100000001000000010000000010000001000000001000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000010000000100000001000000010000000010000000100000001000000100000001000000001000000100000000100000001000000010000000100000001000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000000000000010000001000000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000000100000001000000010000000100000001000000100000001000000010000000100000001000000010000000100000001000000001000000100000010100000100000000100000001100001100100111001011011010000011010110000100110101000000001010110010001100011110,
	960'b000100110001100000100001010000110100110001010100011011001010010011000111010110010000001000000101000000100000011000000100000000110000001100000010000000100000000100000010000000010000000100000001000000010000000100000001000000100000000100000001000000100000001000000001000000100000001000000010000000010000000100000001000000010000000100000001000000010000001000000001000000100000000100000000000000010000000100000001000000100000000100000001000000010000000100000001000000100000001000000001000000010000000100000000000000010000000000000001000000100000000100000010000000010000000100000010000000000000000100000010000000010000000100000001000000000000000100000001000000010000001000000010000000010000001000000001000000010000000100000001000000010000000100000010000000010000000100000010000000010000000100000010000000100000001000000010000000110000001100000010000000010000011000000011000000110000010000000011011101101011110010001111010111110101000000111111001011000001111100011110,
	960'b000101010001101100100011010000000100111001010111011101011010101010111110001110000000001000000100000001000000011000000011000000100000001000000011000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000100000000100000001000000010000001000000001000000010000000100000010000000010000000100000001000000010000001000000001000000010000000100000010000000010000000100000001000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000001000000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000001000000010000000100000001000000010000000010000010100000101000000110000010000000001010101001011110010010111011001100101010001000010001011000001111100011101,
	960'b000100110001110000100101001111110101001001011100011110101010101110110010001000110000001000000100000000110000010000000001000000010000001000000010000000100000000100000010000000010000001000000001000000100000001000000010000000010000001000000001000000010000000100000001000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000000100000001000000010000000100000001000000010000001000000001000000010000001000000001000000010000000000000001000000100000001000000010000000010000000100000001000000010000000100000010000000100000000100000000000000000000000100000001000000100000001000000001000000100000001000000010000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000001000000010000000100000000100000001000000100000010000000100000000010000010000000001001110111011100110011100011011100101010101000110001011000010000100011101,
	960'b000101000001100100100011001111010101010001100001100000011010111010100110000101010000010000000100000000110000010100000010000000110000001000000010000000100000001000000010000000100000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000001000000001000000010000000100000010000000010000001000000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000000100000010000000010000001000000001000000100000000100000001000000010000000100000001000000010000001000000000000000000000001000000010000000100000001000000001000000100000000100000001000000100000000100000001000000100000000100000001000000100000001000000010000000100000001000000010000000100000000100000001000000010000000100000001000000010000000100000010000000010000000100000010000000010000001000000010000000100000001000000001000000100000010000000101000000100000010000000011001011011011010010011111011100100101100001001000001011100010000000011010,
	960'b000101100001110000100011001110110101010101100110100001011010101010011011000100010000010100000100000001000000010100000011000000100000001000000001000000100000000100000010000000010000001000000001000000010000001000000010000000010000000100000001000000010000001000000001000000010000000100000010000000010000001000000010000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000000000000000000000100000001000000010000000100000001000000010000001000000001000000010000000100000010000000010000000100000000000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000000000000010000000100000010000000100000001000000001000000100000001000000001000000100000000100000001000000010000000100000010000000010000000100000010000000100000001000000001000000010000001000000010000000010000001000000010000000010000001100000101000000100000010000000100001001111010111110100000011101110101110001000111001011110010000100011011,
	960'b000100110001100000100100001111010101101001101100100001011010011110011010000101000000010100000011000000110000010100000010000000010000000100000001000000010000001000000001000000100000000100000001000000010000001000000010000000010000000100000000000000010000001000000001000000010000001000000010000000010000001000000010000000100000001000000010000000010000000100000001000000000000000100000010000000010000000100000001000000000000000100000010000000010000001000000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000011000000100000001000000001000000010000001000000010000000100000000100000001000000010000000100000001000000010000001000000001000000010000000100000001000000100000001000000011000000110000001100000011000000010000001100000110000000100000001100000101001010001010111110011111011111000110000101001101001100000010000100011101,
	960'b000100000001101100100100010000100101111001110010100010001010001110100001000110100000010000000100000001000000011100000010000000100000001000000011000000100000001000000001000000100000001000000010000000100000001000000001000000100000000100000001000000010000000100000001000000010000000100000001000000100000001100000010000000100000000100000001000000010000000100000001000000000000000000000001000000010000000100000001000000010000000000000001000000010000000100000010000000000000000000000001000000010000000100000001000000010000000000000001000000100000000100000001000000000000000000000001000000010000000100000001000000000000001000000001000000010000000100000010000000010000000100000010000000010000000100000010000000100000000100000001000000010000000100000001000000010000001000000001000000010000001000000010000000100000001100000011000000010000001100000001000000100000010000000101000000010000010000000101001011111011000010011100100000000110100101010001001100110010000100011100,
	960'b000100100001100100100011010001110110001101111010100100011001111010101001001001000000010000000100000000110000011100000011000000100000000100000010000000100000001000000010000000100000001000000001000000010000000100000001000000100000001000000001000000010000000000000010000000010000000100000001000000100000001000000010000000010000000100000001000000100000000100000001000000010000001000000001000000000000000000000001000000010000000100000001000000010000000100000001000000000000000100000000000000010000000000000001000000010000000100000001000000100000001000000001000000010000000000000000000000010000000100000001000000100000000100000010000000010000000100000010000000100000000100000001000000010000000100000010000000010000000100000001000000010000000100000010000000100000000100000001000000100000001000000010000000100000001000000001000000010000001000000010000000110000010000000101000000110000010000000100001111011011010010011001100001110111000001010110001101100001111100011110,
	960'b000100110001101000100011010010100110100110000010100110101001100010101101001110010000010000000100000000100000010100000011000000110000001000000010000000100000001000000010000000100000001000000010000000010000001000000010000000010000000100000001000000010000000100000010000000010000000100000010000000100000000100000001000000010000001100000010000000010000000100000010000000100000001000000010000000000000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000000000001000000010000000100000010000000100000000100000010000000100000001000000001000000100000001000000010000000110000001000000010000000110000010100000101000000100000011000000011010101001011010110010100100100110111100101011101001101100010000000011101,
	960'b000100100001101000100011010010100111001110001110101010101001010110101110010101010000010000000110000000110000011000000100000000110000001000000010000000100000001000000011000000100000001000000010000000010000000100000010000000100000000100000001000000010000001000000001000000010000001000000001000000010000000100000001000000010000000100000010000000010000000100000001000000100000001000000001000000010000000100000001000000100000001000000010000000010000001000000010000000100000000100000010000000100000001100000010000000010000001000000010000000010000000100000001000000100000000100000001000000010000000100000010000000010000000100000010000000010000000100000001000000100000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000000000001000000001000000100000001000000010000000110000001000000010000000010000000100000010000000110000011000000100000000100000011000000100011100011011000110010110100111111000000001100010001100110010001000011101,
	960'b000100010001101000100001010001010111111010011010101111001001011010101100011101110000100100000110000001000000010000000101000000110000001000000010000000100000001000000010000000010000001000000010000000010000000100000010000000010000000100000001000000010000000100000001000000010000001000000010000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000010000001000000001000000100000000100000001000000100000001000000001000000010000001000000010000000010000001000000010000000100000001000000010000000100000000100000010000000100000000100000001000000010000000100000010000000010000001000000010000000010000000100000001000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000000100000010000000100000001000000010000000100000001000000001000000010000000100000010000000110000011000000010000000110000011000010001100100011010011110011110101011001000101101101010001011010010000000011101,
	960'b000100110001100100100010001110111000100010100101110001111010010110100000100101110001101000000111000001000000001100000111000000110000001000000001000000010000001100000010000000100000000100000010000000010000000100000001000000010000001000000001000000100000000100000010000000100000001000000001000000010000000100000001000000010000000100000001000000010000001000000010000000100000001000000010000000010000001000000010000000100000001000000010000000100000001000000010000000100000001000000001000000010000001000000010000000100000000100000010000000100000001000000010000000100000000100000001000000010000001000000010000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000000000001000000001000000010000000100000010000000100000001000000010000000100000001000000001000000010000001000000011000001000000010100000011000001010000011000101011101010101001100110110011101101101001010001101001001001110010000000011110,
	960'b000100100001101000100000001011101000101010110000110010101100000010010010101010110011111000000101000001010000001100000100000000110000001000000010000000010000001000000001000000100000001000000010000000100000000100000010000000010000000100000001000000100000001000000001000000010000000100000001000000010000001000000001000000010000000100000001000000100000000100000001000000100000001000000010000000100000000100000001000000010000001000000010000000100000001000000010000000100000001000000010000000100000001100000010000000100000001000000010000000100000001000000001000000010000000100000001000000010000000100000010000000100000001000000010000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000100000001000000001000000010000000100000001000000100000001000000010000000100000001100000001000000010000000100000011000001010000001100000100000001110000011101011000101100001001001111001101101111011001111101100000001000110010000100010110,
	960'b000100010001100100100001001000110111011010110111110010101101010110010011101010010111001100001000000001110000001100000011000001010000001000000011000000100000001000000001000000010000001000000010000000100000001000000010000000010000000100000001000000010000000100000001000000100000000100000001000000100000000100000001000000010000000100000001000000100000000100000001000000100000001000000010000000100000000100000000000000000000000100000001000000000000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000001000000001000000010000000100000000000000010000000000000001000000010000000100000001000000010000001000000010000000010000000100000001000000010000000100000001000000100000001000000010000000100000000100000001000000010000001000000001000000100000001000000010000000100000001000000001000000010000000100000011000001010000001000000100000010010001000010001010101001001010000111011000101111001010011001001000001000100010000000011100,
	960'b000101010001011100100000001000000101000110111001110010001101111110101000100110001010000100101001000001100000010000000011000001010000010100000010000000100000001100000010000000100000000100000010000000010000001000000010000000100000001000000010000000100000000100000010000000100000000100000001000000100000001000000001000000010000000100000001000000100000001000000001000000010000001000000010000000100000001000000001000000010000000100000001000000010000000100000010000000100000000100000001000000010000000100000000000000010000001000000010000000010000000100000010000000100000001000000001000000100000000100000001000000000000000100000001000000010000001000000001000000010000000100000001000000010000001000000001000000010000001000000001000000010000000100000001000000010000001000000010000000100000000100000001000000100000001100000001000000100000001000000101000000110000001000000101000001100011110110101001100101001100010011011000101111011010000000101110001001010001111100011001,
	960'b000101100001100100100000001000110010110010100011110000011101011011001110100010111010110001101111000010000000100000000101000000110000011000000011000000100000010000000011000000100000001000000010000000010000000100000010000000100000001000000010000000100000001000000010000000100000000100000001000000010000000100000010000000100000001000000001000000010000000100000000000000000000000100000001000000100000001000000001000000010000001000000011000000100000001000000001000000010000000100000010000000010000001000000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000001000000001000000000000000100000001000000010000000100000010000000100000001000000010000000010000000100000001000000010000000100000010000000010000000100000001000000100000001100000010000000100000001000000000000000010000001000000010000000110000010100000100000000110000010000000110000011100111111010100110100100111101100011001000101101110111101000100010001000110001111100011001,
	960'b000100100001011100011111001001000010000001110001101110111100010011011101101000001001101110100011001011000000010000000110000001000000001100000110000000010000001000000010000000100000001000000010000000100000001000000010000000100000001100000010000000100000000100000010000000100000001000000010000000010000001000000010000000100000000100000010000000100000001000000001000000000000000100000001000000010000000100000001000000010000001000000011000000100000001000000001000000010000001000000010000000100000001000000010000000100000001100000010000000100000001000000010000000010000000100000001000000000000000100000001000000010000001000000010000000100000000000000001000000010000000100000001000000010000000100000001000000100000001000000010000000010000001000000010000000100000001100000010000000010000000100000010000000010000001000000001000000110000010000000010000001000000011100000110010001101010011110010001101101001100101010111001101100010100010000100011001001000010000100011011,
	960'b000100110001101000011110001000100010001000111011101011001011001011001000110001111000100110101000100000010000110100000111000001010000001100000100000001010000001000000010000000010000001000000010000000010000000100000001000000010000000100000010000000010000001000000001000000010000001000000010000000010000000100000010000000110000001000000001000000100000001100000001000000010000000100000001000000010000001000000010000000010000001000000010000000100000001100000010000000100000001000000010000000110000000100000010000000110000001100000010000000100000001000000011000000100000001000000010000000100000001000000011000000100000001000000001000000010000000100000001000000010000000100000000000000010000000100000001000000000000000100000010000000100000001000000001000000100000000100000001000000100000001000000001000000010000001100000100000001110000010000000011000001010000010000011111100101101010001110001111110000011011000010101001100010110010000000100110001001010010000100011100,
	960'b000101010001011100011111001001010010011000100000011110001010001110101010110000111001111110010001101010110101100100000100000001100000001100000100000001010000011000000010000000010000001100000011000000100000000100000001000000010000000100000001000000000000000100000010000000100000000100000001000000010000000100000001000000110000001100000001000000010000001000000001000000010000000100000001000000100000001100000010000000110000001000000011000000100000001100000010000000100000001000000011000000110000001000000011000000010000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000000100000001000000010000000100000010000000010000001000000010000000100000001000000001000000100000000100000001000000010000000100000010000000110000000100000010000000010000000100000010000000010000010000000101000000100000001100000100000001010000101001110001101010101000101110100110101001111001100010100000010010100001111100100110001001000001111100100000,
	960'b000100100001011100011110001000100010010000100101001110101001001010010011101000001011010110001010100111101010010100111111000000110000010100000100000000110000010000000110000001000000001000000011000000100000001000000001000000010000001000000001000000100000000100000010000000100000000100000001000000100000001000000010000000100000001000000011000000100000001000000010000000100000000100000001000000100000001100000001000000100000001000000011000000100000001000000011000000110000001100000011000001000000001100000011000000010000000100000010000000100000001100000011000000110000010000000010000000110000001100000010000000100000001000000010000000010000001000000010000000010000001100000010000000100000001000000010000000100000000100000001000000100000000100000010000000100000000100000010000000100000001000000001000001010000010100000011000001000000010000000101000001100101010110101001100101001000110010010111100010011000101101111001000110110010010100100110001001000010001000011101,
	960'b000100010001100100100001001000010010011000101010001000000101110110001010100010111001011110011100100000101010010110100001001100010000001000000100000001000000001100000011000001100000011000000011000000100000000100000010000000110000001000000010000000110000001100000010000000100000001100000010000000110000010000000001000000010000000100000010000000100000000100000010000000110000001100000010000000110000001100000010000000100000010000000010000000110000010000000010000000100000010000000011000000110000001000000010000000100000001100000011000000110000010000000011000000110000001100000011000000110000001000000010000000100000001000000010000000010000001100000011000000110000001000000010000000110000001000000010000000110000001000000010000000110000001000000010000000100000000100000001000000100000010100000111000001010000001100000011000001000000010000000100010011101010010010011110100000011000100001110110011101001000000100110011000110110010100000100100001000100010001000011111,
	960'b000101010001011100011101001001010010010000100110001000010010101001110101011111011000000010001010100100011000010110100111101000010011011100000010000001000000010100000101000001000000010000000110000001110000010100000010000000100000010000000011000000100000001000000010000000100000000100000001000000100000001100000010000000100000000100000011000000100000001000000010000000110000001000000011000000100000001100000011000000110000001000000010000001000000001100000011000000110000001100000011000000110000001000000011000000110000001100000011000000100000001100000011000000110000001100000010000000110000001100000010000000100000001000000011000000100000001000000010000000110000001000000010000000100000001000000010000000100000001000000010000000100000001000000001000000110000001100000101000001100000011000000011000000110000010100000101000001000000011101010010101001001010000101111110011110110110101101100100011011010101001000011001001010000010100000100111001000110001111000011110,
	960'b000101010001100000011100001000110010001000100110001010000001111100111100011110000111000001110111100000101000010110000101101001101010011001001110000001010000010000000101000001010000010100000011000000110000010100000101000001010000011000000101000001000000010000000011000001010000011000000101000001000000010100000111000001100000010100000101000001000000010100000101000001010000010100000101000001000000010000000100000001000000001100000100000001010000010100000110000001010000010000000101000001010000010000000110000001100000010000000100000001010000010100000101000001010000010000000100000001000000010000000100000001000000010000000100000001000000010100000100000001010000010100000101000001000000010000000100000001000000010000000101000001000000010000000101000001010000010100000011000000100000010000000101000001100000011100000100000100010110011010101000101000100111110001110000011000100101101001011010010110100010000100100001001010000010011100100100001001010010000100011101,
	960'b000100110001100100011110000111110010001100101000001010000010001100011111010011000111000101101110011110000111101110000000100000011010001010110000011110000001110000000000000001010000011000000101000001010000010000000011000000100000010000000011000001000000001100000100000000110000001000000011000000110000010000000100000001000000010000000100000000110000001100000100000001000000001000000011000000110000001100000100000000110000001100000100000000110000010000000011000000110000001100000011000000110000001100000011000000110000001100000100000000100000001100000101000001010000010000000100000000110000010000000101000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000010000000100000000100000001100000100000001000000010100000011000001100000011100000111000001010000010100101100100000111010110010011100011101100110010101100000010110010101000101011001001010110001111100101000001010100010110100100011001000110010001100011101,
	960'b000101010001011000011110000111110010010000100100001010010010100000011100001000000101011001101101011011010111000101110100011111010111111110011000101100001010001001011001000101100000010000000101000010000000011000000101000001000000010100000110000001100000010100000101000001010000010100000100000001010000011000000110000001010000010100000101000001100000010100000101000001000000010100000110000001010000010000000101000001010000011000000101000001010000010100000101000001100000010100000110000001010000011000000101000001010000011000000110000001010000011000000110000001010000010100000101000001010000011100000101000001010000010100000101000001000000010000000101000001100000010100000101000001000000010100000100000001010000011000000100000001010000011100000110000010000000011100000111000010000000010100000100000110100101111010100000101011001001000101110000011000000101100001010111010010110101010000110100000111100010011100101011001010100010101000101000001000010001111100011100,
	960'b000101100001100100011101001000110010001100101000001011010010100000100111000111100010010101010111011011000110100001101110011100111000001010000011100010101010001010110011101000110111001000110101000100000000010000000100000001010000011100001000000010000000100100001000000010000000011100000110000001100000011000000101000001000000011000000101000001100000011000000101000001100000010100000110000001010000010100000110000001110000011100000110000001100000011100000111000010000000011100000111000001110000011100001000000010000000100000000111000010000000011100001001000010010000011100000111000001100000011100000110000001110000011100000110000001010000011000000111000001010000010100000110000001000000010100000101000001100000011100000111000001110000100000001000000001110000011000000110000011110010111001100100100110111010110110011110100000110111000001100001010110000101000101001001010101010011010100100010001001100010100000101011001010110010101100101010001001110010000000011101,
	960'b000100110001011100011110001000100010010100100100001010100010101100101010001001100001110100100001010101110110110001100011011010100110111110000011100100111000101110001101100111111011010010110101100110100111000101010000001110110010111000100101001001000010010000100100001001000010010000100100001000100010000100100001000111110001111100011111001000000010000000100000001000010010000100100010001000100010001100100100001001000010001100100010001000110010001100100011001000110010010000100100001000110010010100100101001000110010010000100100001000100010001000100010001000100010001100100010001000100010001000100010001000100010000100100010001000010010000100100001001000000010001000100011001000000010001000100010001001000010001000100100001001000010011000101011001110010100110101101111100100001010101010101100100111111000100101111110011100010101110101010111010011100100111101011011001101100001111000100101001010000010011100101100001011000010101000100111001000100010000000011101,
	960'b000100010001100100011111001000010010010100101001001001010010110100101101001010000010010000011111001000000100111001101110010111100110000101100110011101001000110010011001100011111000101110010101101000001010110010110010101101011011001110101110101011101011000010110010101101001011011010111001101110101011101110111101101111111011110110111111110000001100000111000010110000111100010011000101110001001100010011000110110001111100011111001000110010001100100011001000110010001100101011001011110010111100101111001010110010101100110011001100110010111100101011001011110010101100100111001001110010001100011111000110110001011100010111000011110000101100000010111110101111001011100110111000101101011011010110110011101100101011000110101110101011001010111010101110101100001011000110101100101000001001001110001000100001011000001001110010010111010101010101001111010101000101110100110011001000000010001100101000001010000010101100100111001011000010101000100010001001010010001100011100,
	960'b000101000001100100011100001001000010001100100110001010010010011100101101001001110010100100100100000111110001110000111101011010110110001101011001011000010110100001110101100010011001001010010101100100111001001010010011100101001001011010011001100110101001110010011101100111111010000010100000101000101010001110100011101001001010001110100100101001101010011110101000101010011010100110101011101010101010101010101100101010111010110110101101101011101010111110110000101100001011000010110000101011111011000010110000101100011011000110110000101100001011000010110001101100001010111110101110101011101010110110101011101010101010100110101000101010001010011010100101101001001010001010011111100111101001111110011110100111011001110110011100100110001001011110010111100101001001000010001101100010101000011110000010011100110110010101011100010100110101000001100000010110010010110000100010001001110010100100101011001010000010101100101011001001100010010100100101001001010001111100011110,
	960'b000101000001011100011100001001000010010000100100001010110010100100101010001011100010100100101000001001010010000000011101001010100101100101101100010110110101011101100011011001010110101101110100100001001001001110010111100101011001010110010100100101001001001110010011100100011000111010001010100001101000010110000011100000111000000110000001100001001000100010001011100011101001001010010110100110001001110010100000101000111010100010101010101011111011000010101111101011111011000110110001101100011011001010101111101011111010110010101101101011101010101010101001101001111010001110011110100110001001010110010001100011101000101010001001100010001000011110000110100001101000011110001000100011011001000010010010100101011001011010010101100101011001011010010110100101101001000010000100011110100110111001100110011000100101111001011011010111110110010001000100001001000010001100100011001001110010100000101100001010100010100000101011001001110010010000101000001000100010000000011111,
	960'b000100100001101000100001001000010010011100101000001001110010100000100111001010010010101100101100001010010010011100100010001000100001111100111000011000110111001001100010010101100101101001100010011001100110110101101111011100000111000101110010011100010111000101110001011011010110101001101000011000110110001101100011011000110110000001011110011000000110001001100101011010110110111001110000011101000111110010000000100001011000100110001011100011101000111110010000100100101001010010010101100101111001100110011000100110001001011110010101100100001000101110001100100010011000000101111101011101110111001101110001011011100110011101100101011000110110001001100001011000010110000101100010011001000110100001101101011100000111010001110101011101100111010101110010011100100110111001101011011001110110001101100010011001010110101101101101010100000010101100100000001000100010010100101001001010100010110100101100001011100010101000101001001010000010011100100010001000100010010100100000,
	960'b000100100001101000011111001000100010010000100110001001100010100000100110001010100010101000101110001010110010101000101001001001010010001100011111001000000100001001110010100011001000000101101011010111000101110101011111011000100110001101101000011011000110110101101010011001100110011001100100011001000110001101100000010111100101101101011010010110110101110001011110011000100110010001100110011001110110110101101111011100100111010101110101011110010111110001111110011111111000000010000001100000011000000110000000100000011000000110000000011111000111100101110110011101000110111001101011011001110110010101100110011001100110010001100011011000010110000101100001011000000101111001011110010111110110000101100001011000010110001101100011011001000110010101100101011001000110010101100110011011000111110110001001011111010101011100101010000111000001111100100100001001010010101100100111001010010010101100101100001010110010100000101010001001100010010000100110001000100010000100011110,
	960'b000101000001011100011100001001010010010000100100001010010010100000101000001010100010110000101001001011000010111000100111001010000010100000100101000111110001111000100101010011001000011010101111101100111010011010011011100110011001101110011100100111001001110010011100100110111001110010011100100110101001100110010111100101101001001110010011100101001001001110010100100101011001010110010101100101111001011110011000100110101001101010011010100111111010000010100000101000101010001110100011101000111010010010100100101000111010001010100001100111111001111010011011100110111001011010010101100101001001000110010001100100001001000010001111100011101000111010010000100100001000111010001101100011111000111110010001100100011001001010010001100100111001001110010001100100101001101110100111101000111000001101010011001010110001101100011111001001110010100000101001001010000010011100101100001010000010100100101110001010000010100100101100001001100010010000100101001001000001110000011111,
	960'b000101000001101000011101001000010010000100100110001010000010011100101100001010000010110000101011001010100010110100101001001010100010101000101000001001100010000100011111000111000001110100110110010111010111100010000101100001111000100010001000100010011000100110001010100011001000100110001011100011001000110010001011100010101000100010000111100001011000100010001001100010011000101010001100100011101000111110001101100011101001001110010101100101111001100110011100100111101010000010100000100111101010001010100011101000011010000010011110100110111001100010010100100011001000111010001110100010111000100110000111100001101000010010000101100000101000010010000110100001111000100010001010100010011000101110001001100011001000101110001010100010101000011110000111100001100111100001011011001110100010010000011111001000110010100100101010001011010010110000101001001010100010100100101010001010110010100000101000001010010010110100101001001010100010100000100100001000110010000000011011,
	960'b000100100001100000011110000111110010010000100110001001100010110100101110001011000010100000101100001010110010011100101011001010100010011100101010001010110010101100101001001010000010010100100010000111100010000100100100001011110101000000110010001000110010000100100111010010110100000000101011001001100010011000100100001000010010100101010001001111010010010100100010001000110010010000100100001000110010101101010001001111110010101000100101001001000010001100100100001001000010100101010000010000100010101000100101001001110010011100100110001001000010011101001001010010000010101000100011001001000010010000100010001000100010010001000111010011000010101000100010001000100010000100100010001001010100111000111111001010000010001100100010001110110100110100101011001000100001111100011110001000010010011000101010001011110010110000101100001001110010100000101110001011100010110000100111001010010010110000100111001011000010101100101001001011000010101100100100000111110001111100011101,
	960'b000110000001100000011010001000000010001100100011001010100010101000101101001011010010110000101000001010010010100100100111001010100010111000101011001010110010100000101010001010010010100000101000001001110010011100101001001100100100011001000011001010000010011100101100001110100100110100101110001001010010011000100111001001010010101000111101010001110010101000100101001001010010010000100100001000100010011100111001010001110010011100100011001000000001111100100001001000000010001000111000010010100010010000011101000111010001111000011110000111100010010100110100010010010010110100100010001000010010000100100000001000010010010100110101010011000011001000100101001001010010010000100101001010010011101001001100001010110010011000101000001101000100110100110111001010110010101100101101001011110010111000101111001010100010100100101000001010100010111100101100001011010010110000101111001010110010100000101001001010000010101100101111001010100010100100101000001001000001111000011100,
	960'b000110000001101000011011001000000010000100100110001010100010100100101100001011000010111000101010001010010010101000101010001011000011001000101010001011010010110100101110001010000010011000100111001010000010101100101100001011010011000000110000001011010010111000101101001011010010110000101110001010110010111000101100001011010010101000101110001100000010110100101101001011100010110000101100001011000010110000101100001010100010100100101000001010010010101100101010001010010010101000101100001011000010100000100111001001110010100000101010001010000010101000101100001010110010101000101000001010010010101000101011001011010010110000101111001100010010110100101101001011010010101100101011001011000010111000101111001011010010101100101101001011100011000000101110001011110010101100101100001010110010101000100111001010100010100100101001001010000010111000101011001011000010101100101110001010110010101000101001001010100010101000101101001010100010100100101000001000110001111100011101,
	960'b000100100001100000011101000111010010001100100101001001110010111000101100001010110010100100101010001010110010101100101101001010010010101000110000001011100010110100101010001010110010101000101010001010010010010100101000001010110010101100101000001010000010100100100111001010000010011100100111001010010010101000101000001001110010100100101010001010010010011100101000001010000010101000101001001010110010011100100110001010010010011100101001001010010010100000101010001010010010100100100111001010000010100100100111001010000010100000100111001010100010101000101000001001110010011100100111001010000010100100100101001010000010101100101010001001100010100100100110001001000010100100101001001001100010101000101001001001110010100000101000001001100010100000101001001010000010100100101011001011010010100100101100001011010010101100101100001010100010100000101111001011100010110000101001001010110010100100101001001011000010101000101000001100000010101100100101001000100010001100011110,
	960'b000100110001101000011100000111110010001100100110001001110010100100101110001010010010101100101101001010010010101000101011001011010010100100101111001011110010100000101100001011100010101100101010001011010010101000100111001011010010110000101011001011000010101100101001001010110010101100101010001010000010111000101011001010110010101100101010001011000010110000101101001010010010101000101110001010010010101100101101001010110010101000101011001011000010100000101101001011110010101000101100001011000010101000101001001010110010110000101001001010110010110000101001001011000010101000101001001010000010101100101011001010010010110000101010001010100010101100101000001001110010100100101101001010100010101100101010001010100010101100101010001011010010110000101100001011000010101000110000001010010010101100101110001010100010101000101001001011010010110000101001001011010010101000101101001010110010101000101011001010110010110100101011001010010010100000100011001001100010000100011100,
	960'b000101010001011000011011001000110010000000100011001010010010100000101011001010110010110000101001001011010010111100101010001010110010110000101010001010110010101100101101001010100010111100101110001010100010110000101011001010110010101000101011001010100010100000101111001011010010100100101100001010100010101100101001001011100010100100101011001011110010101100101001001011010010100100101101001010100010110100101010001011000010111000101000001010110010110000101001001010100010101000101101001010000010110000101111001010010010101100101101001011000010101100101011001010110010100100101111001011010010100000101100001010100010100100100110001010110010100100101100001011000010010000101010001010100010100100101010001010110010100100101010001100000010111000101000001010110010101100101011001010110010110000101000001010110011000000101011001010100010111000101010001010110010101100101101001010000010101100110001001010110010101000101100001010000010011000100110001001000001111100100000,
	960'b000100110001011000011011001000000010000000100101001010000010100000101000001011000010101000101100001010110010110000101011001010110010110100101000001001110010110100101001001010010010110100101110001010110010101100101100001010010010100100101011001010010010101000101101001010110010101000101010001011000010100000101011001011000010101000101011001011000010101000101001001010110010101000101000001011100010101000101000001010110010111100101010001010010010101100101000001001100010101100101010001010110010110000101101001011000010101100101101001010100010100100101101001010100010101100101011001010100010100100101001001011000010011100100111001011000010100100101000001010010010100100101001001010100010011100101001001010100010101100101101001011100010101100101100001010110010101100100110001010100010101000101001001010110010110100101100001011000010101100101001001001110010101000101001001010100010101000101101001011010010101000101001001010000010010100100110001000010010000100011100,
	960'b000100110001101100100000000111110010011100101001001001000010011000101011001010100010101100110000001011100010101100101110001011000010100000101000001010100010100100101010001011110010110000101011001100100010110100101001001010100010101100101000001011010011000000101100001011110011000000101010001010000010101100101001001010000010110000101110001010010011000000101110001010110010100100101011001010010010100100101110001011000010101000110010001010110010011100101000001011010010100100101011001100100010111000101100001100000010101100101000001010010010101100100110001010010011000000101011001011000010111100101001001001100010100000101000001010000010110100101001001010100010111000101011001001110010101000101010001010000010110000101110001011000010110100101111001011000010100000101001001010010010100100101100001011110010101000101110001011110010100100100111001010110010100100101000001011100010111000101100001100010010110100100110001001110010011100100011001000100010001100011101,
	960'b000100110001011100011011001000010010001000100101001001010010100000101001001011000010101000101001001010100010111000101010001010100010101100100111001010000010110100101001001010110010110000101100001011000010100100101100001010100010100100101100001010100010101100101100001010110010101000101001001010100010100000101011001010100010101000101100001011100010101000101011001010110010101100101001001011010010101000101001001010100010110000101010001010000010110000101000001001110010101100101011001010110010100100101101001010010010100100101011001010100010100100101100001001110010100000101101001010100010011000100111001010100010011100101001001011000010100000101011001011000010011100101000001010110010100000101010001011010010101000101001001100000010110000101001001011000010101100101000001011000010101100101000001010010010111100101011001010100010110000101100001010010010101100101011001010100010110100101111001010010010100000101011001010000010011000100110001000100001111100011110,
	960'b000101010001011100011010001000100010000000100011001001100010010000100110001001110010110000100111001010110010111000100111001010100010100000100101001001110010100000101010001010000010110000101100001001110010101100101001001010010010011100101010001010110010011100101100001010110010011000101010001001100010100100100110001011000010100000101000001011100010100000101001001011000010011000101001001001100010101100100111001010100010111000100111001010000010100100100111001001110010011100101100001001100010100100101011001001100010100100101001001010010010100000101001001010110010011000101100001010010010010000101011001001010010011100100100001010010010011000101001001010100010010000101010001001110010011100100101001011000010101100101000001011010010100000101000001010110010011000101011001001110010101100101001001001110010110000101000001010100010110000101000001010110010011100101101001010100010100100101100001001110010101100101001001001100010011000100100001000110001110100011101,
	960'b000100100001100100011100000111100010000000100110001000110010011000101001001001100010011000101001001001100010011000101001001010000010010100101000001010010010010100101000001010110010011100100110001010100010100100100111001010110010101000100110001010010010100000100111001001110010100100100111001001010010110000101001001001100010101000100111001001010010100000101001001001100010101000101100001001010010011000101001001001100010011000101001001010000010010100101011001010100010010100100110001010010010011100100101001010100010100100100110001010110010101100100110001010100010100000100110001001000010100000100101001001010010101000100111001001010010101000100110001001100010100100100110001001010010110000101010001001010010100100101000001001010010100000101001001001010010100000101010001010000010010100101001001010000010010100101000001010010010010000101011001011000010100100100101001010100010100000100101001010100010100100100011001010010010100000100011001000010001111100011010,
	960'b000100000001010100011011000111000010000000100001001001010010011100101000001001110010001100100101001001010010010000100101001000110010011000100111001010000010011000100001001001010010011000100110001001010010010000100111001010010010100000100111001000110010011000100111001001110010001100100100001001100010100000101000001001010010010100100101001001000010011100100001001001010010101000101001001001110010001000100100001001100010001100100111001000110010011100101001001010010010100000100010001001000010011000100100001001000010010000100101001010000010100000100111001000110010001100100011001001010010001000100010001001100010011100100110001001100010011100100110001001100010010000100100001001110010100000101000001001100010001100100110001001000010011000100011001001100010011000100111001001100010011000100010001001100010001100100110001000100010011000101000001010000010100100100101001001000010011000100110001001010010001000100110001001010010010100100011000111110001110000011000,
	960'b000100010001010000010111000111000001110000100010001001010010001100100111001001000010011100100011001000100010001100100010001001010010011100100101001001010010010100100101001000010010001000100010001000110010011100100101001001100010001100100110001001100010010000100100001000100010010100100111001001000010001100100011001010010010011100100010001000110010001000100100001001100010010100100101001001010010100000100101001000100010001100100011001001110010011100100100001001000010001100100111001001000010010000100011001000110010011100101000001001000010001100100101001001010010000100100010001000000010001100100101001000110010001100100100001001110010001100100011001000100010001000101000001001100010010000100011001001100010010100100010001001000010001100100111001001110010010000100100001001000010011000100110001000110010010100100010001001100010100000100011001001010010010000101000001001010010001100100100001001000010011100100111001000110010001000100010001000100001101100010110,
	960'b000011110000111100010101000110000001101100011101001000100010000100100010001000100010001000100000001000010010000000100000000111110010001000100001001000010010001000100000000111100010000000100000000111110010000000100010001000100010000100100011000111110010000000100000001000000001111100100001001000100010001100100010001000110001111000100000001000000010000100011111001001000010001100100011001000100010001000100000000111110010000000100000001000000010001100100010001000110010001000100001000111110010000100011101000111110001111000100011001000100010000000100011000111110001111100100000000111100001111000011111001000010010000100100000001000100010000000100000001000000001111100100000001000100010001000100010001000100001111100100010001000010010000100011111001000010010001000100010001000100010000100011110000111110010000000100001000111110010000100100011001000100010000100100000001000000010001000100000001000010001111000100001001000010010000000011110000110100001100000010111,
	960'b000011100001000100010101000101110001101000011011000110100010000000011111000111000001101100011111001000000001111000011111000111010001110100100001001000000001101100011101000111110001111000011111001000010001110000011101001000100010000100011100000111110010000000011011000111100001111100011011000111100010001100100010000110110001111100100000000111000010000100011111000111010010000100100010000111110001110000011110000111010001110000011111000111000001101100100001001000010001111000011101001000010001111100011011000111110001110100011011001000100010001000011100000111100010000000011100000111010010000000011011000111010010000100011111000110110010000000011101000111110001111100011100000111010010000100011111000110100010000100100001000111010001111100011110000110110001111000100001000111100001101100011111000111010001101000011110000111100001101000100001001000010001110100011100001000100001111100011100000111100001111000011011001000010010000000011001000110100001100000010011,
};
localparam [0:85][959:0] g_picture = {
	960'b000011010000110100001110000100000001001000010010000101000001011100010111000101110001011000010101000101100001010100010111000101010001011100011000000101110001011000010101000101010001011000010101000101100001010100010110000101110001011100010111000101010001011000010110000101010001010100010101000101100001011100010111000101100001010100010101000101010001010100010100000101000001011000010110000101100001010100010100000101100001010000010110000101000001011000010111000101110001010100010100000101010001011000010101000101100001010000010110000110000001100000010110000101000001010100010101000101010001010000010010000101000001011000010110000101010001011000010110000101010001011000010101000101000001100100011001000101100001011000010110000101010001011000010110000101100001011100011000000101110001010100010101000101100001010100010110000101010001010000010111000101110001011100010100000101010001011000010101000101110001010100010100000101110001010100010011000100000001000100001110,
	960'b000011010000111100010010000100110001011100011010000110010001101100011110000111000001101100011110000111000001101000011100000111100001101100011101000111100001101100011011000111010001110000011010000111000001101100011001000111010001110100011010000111000001110100011010000110100001110000011011000110100001111000011110000110110001110000011100000110100001110000011101000110100001101100011110000111000001100100011011000110100001100100011011000110110001100000011011000110110001101000011010000111000001100000010111000110110001110000011010000111000001110100011011000110110001101100011000000101110001101100011010000110000001110100011100000110100001110000011011000110100001110000011101000110110001110100011110000110110001110100011100000110110001101000011100000111010001101100011111000111000001101000011101000111000001101100011011000111000001101100011010000111000001101100011010000111000001101100011010000110110001110000011011000110100001101100010111000101010001010000010001,
	960'b000011110001001100010100000110100001101100011100001000000001111100100001000111110010001100100000001000000010001100100001001000000010001100011111001000110001111000100010001000000010000100100011001000000010000100100010001000000010000100011111001000100001111100100001001000010001111100100010001000010010000000011111001000000010000000011111001000010010000000100001001000010001111000100001000111110010001000100000000111110010001000011110001000000010000100011101000111110001111100100010000111110001111000011111000111010010000000100001000111100001111000011110001000010001111000011110000111100001110100100000000111100010000000011110000111110010000000100001001000110001111000100000001000100010000000100000001000100010000100011111001000100010001100100000001000010010000100100001000111110010001000100000000111110010010100100010001000000010001100100001001000010001111100100010000111110010000000100011001000000001111100100010000111100001111000011011000110110001011000010100,
	960'b000100010001010100011001001000000001111100100000001000110010010000100010001001010010011000100100001001100010100100100111001001000010010100100101001000110010011100100110001001000010011100101001001001010010010100101000001001010010010000100111001001010010010000101000001010000010010000100100001001110010001100100101001010000010010100100101001010010010011100100100001001010010010100100011001001010010011000100100001001000010100100100101001000110010011000100100001000010010010000100100001000110010011000101010001000110010001100100111001001000010001100100111001001000010010100100110001001110010010000100010001001000010000100100000001000110010010000100110001001110010010100100100001001100010010000100100001001100010011000100111001010000010100000101000001001010010011000100011001000110010011000100101001001100010101000100111001001110010011000100110001000110010010100100101001001000010011000101010001001010010010100100101001001000010000000100010000111110001110100011001,
	960'b000100010001100000011111001000010010011000101001001001100010011000101011001010100010101000101101001011110010110000101111001011100010100100101000001010100010100000101010001011100010101100101100001100000010110000101000001010010010101000100111001010010010111100101011001010110010111100101001001001110010101000101010001010010010101100101111001011000010111000101110001010000010100000101010001010000010011000101101001010110010101000101110001011000010010100100111001010010010011000100111001011010010110000101011001010110010101000101000001010010010100100101000001010010010111000101100001011010010111100101001001001010010011100100110001000110010101100101100001010110010111000101011001001110010101000101011001010010010110000101110001011000010110100110000001010110010100000101001001010010010100000101100001011100010110000101110001011110010100100101000001010110010011100101000001011010010111000101011001011100010110100100111001001110010100100100011001000000010001000011101,
	960'b000101000001011100011110001001000010011100101001001010100010110000101100001011110010111000101110001011110011001000101111001011110010111100101100001011000010111100101101001011110010111100110001001100000010110100101101001010110010110100101111001011010010111000101110001011100010111100101100001011010010101100101101001011010010101100101110001100010011000000110000001011000010111000101101001011110010110000101111001011110011000000101110001011100010110000101011001010110010110100101101001011110010110100101111001011010010110000101110001010110010101100101110001011010010110100101110001100000010110100101011001011010010101100101011001011000010101000110000001100000010101100101100001100000010110000101100001100000010110100101110001100010011000000101110001011010010111100101100001011000010111000101101001011100011000100101111001011010010110100101111001011100010111100101111001011010010111000110001001011010010110000101110001010110010100000101001001000110010000000011110,
	960'b000110000001101000100000001010010010011100101000001100000010111000110000001011110011001100101111001100010011011100110001001100100011010100101111001100100011000000110010001011010011000100110101001011110011000000110001001011100011000000110011001100110010111000110100001101000010111000110001001011110010111100110000001100110011000000101111001101110011001000101111001100110010111000101111001100000011001100101110001100010011011000101110001011110011001100101100001011100010111000110010001011010011000100110101001011110011000000110000001011100010111100110001001100010010110000110100001101010010110100110001001011110010111100101111001011110010111000110010001101000010111000110001001100100011000000101110001100010011001100110000001101010011010000110001001101010011000100110001001011110011000100110010001011100011010000110001001011110011010000101111001100100010111100110100001100010011000000110101001100010011000000110010001010110010110100101001001010010010000100100000,
	960'b000101110001111000100001001001110010100100110000001100010011000100111000001100100011010000110110001100100011001100110011001101110011010000110100001110000011001100110101001101000011001000110010001100110011011000110011001101100011011100110010001101100011010100110010001100110011010100110110001100010011011100110101001101000011011100110010001100100011000000110101001101010011001000110111001100110011001100110100001100010011001000110010001101010011001100110010001101100011000000110011001100100010111100110001001100100011010100110001001100110011011000110001001100100011001000110001001100010011001100110100001011110011010100110110001011110011011000110010001100100011010100110110001100010011100100110111001100010011010100110110001100100011001000111000001101010011001000110111001101110011001000110101001100110011000100110010001101100011010000110101001110010011010000110011001101100011001100110011001101000011011000110010001100110011010000101101001010010010011100100001,
	960'b000101100001110100100100001001110010110000110001001100010011011000111010001110100011001000110101001101110011001100111001001101110011001000111000001101110011011100110100001101010011011100110010001101110011010100110100001111010011110000110101001101000011011100110101001101000011100000110101001101010011101100111010001100010011010000110110001100010011011000110101001100100011100000111011001110000011001000110101001101100011001000110111001101010011000100111001001110010011010100110010001101000011010000110001001101010011001100110011001110010011101100110100001100100011011100110100001100100011011000110011001100110011100100111000001100010011010100110101001101010011100000110101001101110011100100111010001101100011001000110101001100100011010100110110001101000011010100110101001101100011011100110010001101100011001100110101001101000011010000111000001110100011011100110100001101000011011100110011001101100011010000110100001101110011010000101110001010000010011000100001,
	960'b000110110001111100100011001010100010110000110001001110100011011100111001001110100011101100110101001101000011011100110110001110100011110100111000001101110011101000111011001101000011010000110110001100110011100000111110001110010011100000111010001110010011011000110110001101100011010100111001001111000011100100111000001110100011011000110011001101000011010000110100001110110011100000110111001101110011101100110111001101000011011000110011001101000011110000110111001110000011100100111011001101010011001100110101001101000011011000111101001101010011011100111100001110010011001100110011001101000011010000111000001110000011100000110100001110000011011000110110001110000011011000111011001111100011100000111001001110110011101000110101001101100011010000111001001111100011101100110111001101110011110100111011001101000011011100110100001101110011110100111011001110010011100100111101001110000011001100110111001100110011011100111101001101010011010000110010001011110010011100100000,
	960'b000111000010000000100100001010010010110100110000001110000011011100111010001110010011101000110101001101000011011000110110001101010011110100111000001110010011101000111010001101010011010100110100001101000011011100111101001110000011100000111001001110010011010100110101001101010011010000111000001111000011100000110110001110100011010100110011001101000011010000110100001110100011100000111000001101100011101000110110001100100011001100110001001101010011110100110111001110000011100100111010001101000011010100110110001101010011010000111010001101100011011100111001001101010011001100110011001101000011001000110111001110000011100100110110001101100011011000110110001101100011011100110101001110110011100000111001001110010011010100110100001100110011010100110100001101110011101000111001001110010011101000110101001101100011010100110011001101000011100000111010001110100011011100111001001100110011011000110101001101100011010000111011001101100011010000110000001010110010011000100010,
	960'b000110000010000000100110001010010011000000110010001100100011101000111101001110100011010100111000001110010011010100111001001110010011010000111100001111000011100100110101001110100011100100110101001110100011100000111010010000110100001100111110001111000011111100111101001111100100000000111101010000000100011001000100001111010011111001000000001111000011111000111110001110010100001001000100010000100011110100111111010000000011101100111110001111100011110101000101010000110100001000111011001111110011111100111101010000000011110100111010010001000100001100111101001111000100000000111110001111100011111100111100001111000100001101000011001110110100000000111111001111100100010001000001001111000100010101000101001111010011111101000000001111010011111001000001001111010011100100111111001111010011001100111010001110110011010100111000001110100011010100111010001111010011110000110010001110000011101000110011001110010011101100110100001110100011101000110000001010100010100100100011,
	960'b000110010010000000100101001010100010110100110101001101110011010100111011001101100011010100110101001101100011101100110110001110110011100100110110001111000011010000111010001111010011101101000100010011000101100101100000011010100111000001101110011100010111000101101101011011010111000001101111011010110110111001101101011011000110111001101101011011100110110001101110011011000110110001110000011010010110100101101100011010000110011101100110011010100110100001101000011010100110010101101000011010000110010101100110011001100110101001100111011010000110101001101000011010100110100001101010011011000110110001101110011010100110110101101011011010100110110001101101011011010110110001110000011011100110111001101111011011100110110101101101011100100111000001101011011010010101101101010100010001100100000101000000001101110011100100110111001110000011101100110101001110110011010100111001001110010011010100111000001101100011101000111001001100100011001100101111001011100010011100100011,
	960'b000110100001110100100100001011110010111100101111001101100011011100110110001110000011011100110010001110000100000000111000001101110011101000110111001110010011110001001010010100000110101010000111100101001001001010000011011110100111100101110100011011010110100001100100010111110101100101010100010011100100110101001100010010110100101101001011010011000100111001001011010011000100101101010001101000011010110110101100101100101011110111000010110001111100110011010000110100111101001011010100110100101101001011010011110011111100110011001000110000011011101110110010101010111010110010011001010011100100101001001010010010010100101101001100010011000100110001001101010011110100111001001110010100000101010101011011011000010110010001101000011100000111101001111011011111011000011010010011100100000111111001100001010011000100100000111111001101100011101000111000001101100011011100111010001101010011100000111110001101110011010000111010001101010011000000110010001011010010011000100100,
	960'b000110000001111100100110001011010010111100110010001100100011010100110011001101110011011000111001001110110011101100111100001110100011100000111100010001100110000110000111101001011001110001110101010011110011001000101010001001100010100000100111001010010010101000101010001010110010100100101001001010100010100100101000001001110010010100100101001000110010001100100011001001010010010100100011010100001010100110110101101111001100010111010010110111011110011111101100111100101111010111110110111101101111010111110011111011011110011111011110110101011100011010111100101101111010001001000110001000110010010100100101001001110010100000101001001001110010100000101010001010100010101000101001001010100010101000101100001010100010101100101010001011010010111100101110001011010011000000111101010110001000000110011110100111010111101001011001010010110011101000110111001101010011010100110110001110100011101000111000001110110011101000110110001100110011000100101111001010110010110000100101,
	960'b000101110001111100101000001010110011000100110110001100010011001000111000001101110011010100111010001110110011101100111101010000000100011001100010100100101010011010000010010011010010110100101000001011010011001000110101001100100011001000110010001100010011000000110001001011110010111000101110001011100010110000101101001011010010110100101101001010110010101100101011001011010010111000101101001001010011100001101110100011111001100010011101101000001010001110100101101001111010100010101001101010001010100010100111101001101010010010100001100111011001100010001111011011000011011000100110001010110010101100101100001011000010101100101011001010110010101100101101001011100010111000101110001011100011000100110100001101100011101000111010001111000011101000111010001110100011100100111001001101000011000000110100010101101000100010100010100001010101011101000010001110010011010100110101001110000011101000111001001110110011101000110101001100110011001100110000001010110010101000100100,
	960'b000110100001111000100100001011110010111000101111001101010011011100110110001110000011110000111000001110100100000101000010010101111000100110100010011011100011011100101011001100000011011100111010001110100011011100110101001101100011011100111010001110010011101000111001001110010011100100111001001101110011011100110111001101110011100000110110001101110011100000111000001110000011100000110111001110000011010100110000001100010011001100110011001100100011001100110010001100010011000000101111001011110011000000110000001100000011000000110000001100100011000100110001001100100011011000110110001101010011010100110101001101000011010100110101001110000011100000111001001110100011101100111010001110110011101100111010001110110011110000111100010000000100001101000001010000100011111101000000001111110011110100111011001101010010110001000010011110111001110101110110010011100011111000111100001101110011011100111110001101100011001100111001001101000011000100110001001011010010011000100100,
	960'b000110010001111100100100001010110010101100110001001110010011010100111000001101010011110000111001001110100100110001101011100111010111100000110101001010000011001000110111001110110011111101001000010111000111001110000111100101001001111010100000101000001010000010100001101000011010000110100001101000101010001110100100101001001010010110100101101001111010100010101001101010011010100110101010101010011010101010101010101010011010100110101001101010011010100110101010101010011010100110101001101010011010100110101001101010011010100010101000101010011010100110101001101010001010100010100111101001111010011010100101101000111010010010100011101000111010001010100010101000011010000110100001101000111010001110100100101001011010011110100111101010001010100010100101100110101000101101110101011000000100101101000000001110110011101000110100001010010100001010000110100011010101101001000011001110110011011100111001001101100011101000111001001100110011010100101111001011100010100100100011,
	960'b000101100010000000100110001010010010111100110110001100110011100000111110001110100011010101000000010011100111101010010010010011100010110100110101001110010011101101000101011000101000101010101101110000111100110111001011110001001011110110111010101101111011011010110111101101101011011010110100101101001011010110110101101101011011011010110111101101101011011110110111101110011011101010111010101110111011101110111100101110111011110010111011101111001011110010111100101111001011110010111100101111001011110010111011101111001011110010111100101111011011110110111110101111101011111010111110101111101011111010111110101111101011110010111100101111001011101110111011101110111011101010111011101110111011110010111101101111101011111110111111101111111100000111000100110011001101001011010000110000111010011110000011010111000100010100111100001101110011001100101110010111011001000001100111010001100011101100110101001110100011101000110011001110010011101100110001001010110010100100100100,
	960'b000110110001101100100100001010000010111100110001001101010011100000111011001110110011110101001100100001100111111100111111001111000100001101000110010010100110101010011101110000111101000011000011101000111000000001100111010110000101000001001110010011010100110101001110010011100100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001110010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110001001100010011010100110101001101010011010100110101001110010011100100111001001111010011100100111001001110010011100100111001001110010011100100111101001110010011100100111001001110010011110100111101001110010011100100110101001101010011100100111001010001010110100110101010000110101010001100011011001101101110001001000001011111010001110100001001000000001101010100100110000011011100000100011100111010001101110011011000111011001101110011011000110100001011010010011000100010,
	960'b000111000001111100100011001010100010101000110011001110100011100100111011001111110101011010000110011100100100000101001011010100000101101101100110100101011100001011001110101100010111100101010010010001010100100101010010010111010110001101100101011001110110011101100101011001000110001101100011011000100110000101011111010111110101111001011110010111100101110101011101010111010101110101011101010111000101110101011110010111100110000001100000011000000110000101100010011000110110001101100101011001010110010101100101011001010110010001100011011000110110001001100000011000000101111101011110010111100101110101011101010111010101110101011101010111010101110101011101010111010101111001011111010111110110000001100001011000100110001101100100011001010110011001100010010110110101000101000111010001010101011010000010101101101100101110110101100000100101100001010011010011110100001000111111011110110111000101001000001101100011100100111110001101110011011100110101001100000010100000100011,
	960'b000110010001110100100101001010000010111000110000001101010011101101000000010100001000001101101110010010010101100001100101011100110111110110110000110011001011011101110010010001110100101001011110011100011000001110001101100100111001011110011010100110001001100010010101100101001001001010010000100011101000110110001010100010001000011010000101100001001000001110000010100000011000001110000100100000111000010010000100100001101000100010001001100011001000110110010000100100001001001110010110100101111001011110010110100101101001010110010011100100001000111010001100100010111000100010000110100001101000010110000100100001001000001010000010100000111000010010000100100001011000011010001000100010101000110010001101100011111001001010010100100101101001011110010110100101011000111010000100011100000101101001001000010011000111110110111100110000111001110101101000011000000110000001010011010000100111100001101100010001100011011100110111001110110011100100110010001011000010100000100100,
	960'b000101100010000000100101001010000010111100110101001100100011101001001111011110010111001101001000011000000111100110000111100011001011101111001011100100100100110101001101011001100111111010001001100011011000111010001101100011001000101110001100100010101000101110001010100010101000100010000111100001001000001110000001011111111000000001111111011111010111110101111101011111010111110101111101011110110111110001111101011111100111111110000000100000111000001110000110100001111000100010001001100010101000100110001010100010101000100110001000100001101000010110000011100000011000000001111111011111100111110101111100011111010111101101111011011111000111110001111100011111010111111101111111100000101000001010000100100001011000011110001001100010101000101110001100100011101001000010010100100101001001000110000000011001010100101101010011100111101100010010100111011100110110110101101100010101110100010001110111011001110100010000110100001101100011011100101110001011100010101000100010,
	960'b000110100001111100100100001011010010111000110001001101110011111001101111011111010100101001011101100000011001001110010011110000001100001001110000010001110110010110000011100010111000101010000110100000111000010010001001100011011000111110010001100100001001000110010000100100001000111110001110100011001000101110001001100010011000100110001000100001111000011110001000100010001000100010001000100001101000011110001000100001111000100110001001100010101000101110001110100011101000111010001110100011111000111110010000100011111000111110001110100011011000110110001010100010011000100110001000100010001000011110000111100001111000011110000111100001101000011010000110100001101000100010001000100010011000101010001011100011001000111010010000100011111000111110010000100011011000100110000110100001111000101010010000100100001000000101011110010001111000000011000000101010010111011101111010011010000101001101000110011110100101110000111111001100100011000000110000001011100010010000100100,
	960'b000110100001111000100100001011010010111100101111001110010101110010000011010010110101011101111001100011001000111110111111101111010110000101010001011111001001000010001100100001001000000110000100100011111001001010010001100011011000101010001001100001111000011110000110100001101000011010000110100001001000001110000010100000111000001010000010100000011000000110000000100000001000000110000000100000011000000110000001100000011000000110000010100000111000001110000101100001011000011010000101100001111000011110000111100001101000010110000101100001001000001010000010100000111000001110000010100000101000001010000001100000001000000010000001100000001000000110000001100000011000000110000001100000111000001110000101100001101000011010000110100001111000101010001101100100011001010010010011100011001000001110000010100010001001000010010011011101010100101101110000101110101010001101111000011110110110000101000111010010110111100001001110001101010010111100110010001010110010100000100100,
	960'b000110000010000000101000001010110011001000110101010001110111111101010011010010100110011110000101100000111011101010111101010111110101100110001101100101111000101110000100100001001000111110010001100010000111111001111100011111000111110001111100011111000111110001111011011110110111101001111010011110010111100001111000011101110111011001110110011101110111011001110110011101100111011001110110011101100111011001110110011101110111100001111000011110000111100001111001011110010111101001111010011110100111101001111010011110100111101001111010011110000111011101110111011110000111100001110111011101110111011101110110011101100111011001110111011101100111011101110110011101100111011001110111011101110111011101111001011110010111101001111010011110110111110001111100011110110111110010000010100011001001010010001110100001001000100010010000100110111000100001010010011011101011011110011001011100110110111101010011001101100101101001101100001111100011001100101110001010100010110100100111,
	960'b000110000001111100100101001011000010111000111011011010100110111100110110010011110111000101111011101100011100001001100110010111011001011010011010100011111000011110001111100101001000010101111011011110010111101001111011011110110111101001111011011110110111101101111011011110110111101001111010011110010111100001111000011101110111011001110110011101100111011101110111011101100111011101111000011110000111011101110111011110000111011101111000011110000111100001111001011110010111100001111001011110010111100101111010011110100111101101111010011110000111100001111000011101110111011101110111011101110111011101110110011101100111100001111001011110010111011001110111011101110111100001110111011110000111100101111001011110010111100101111001011110100111101001111011011110110111110001111100011110110111111110001101100101011000101010001000100100111001110110010100010101100111100010110010100010010110011101011100010000010010111001110001010101010011001100110010001011000010011100100100,
	960'b000110100001111000100011001011010010111101001001100000110011101100111001010110000110011010100001110001010111110101011011100111001001110110010001100010111001011010010001011111010111100101111011011110010111100101111001011110010111100001111001011110010111100101111000011110000111100101111001011110000111100001111000011110000111011101110111011101100111011101110111011101100111100001111000011110000111100001111000011101110111100001111000011101110111011101110111011110000111100001111000011110000111100001111010011110100111100101111000011110000111100001111000011110000111100001110111011110000111100001111000011110000111100001110111011110000111100001110111011101100111011001110110011110000111011101111000011101110111100001111001011110010111100101111001011110010111101001111011011111000111110101111101100001101001101010010011100011011001011110100100100101110101010110001100101001110111010101011000010001000010101101000001011100010011110100101101001011100010010100100011,
	960'b000110000010000000100011001010000011010001101100011000110010110000111100010100101000001011000000101000000101011010011000101000101001010110001101100110011000111101111110011110110111101001111011011110010111100001111000011110000111100001111000011110000111100001111001011110000111100001111000011110000111011101110110011101110111100001110111011110000111100001111000011110000111011101110111011110000111100001111000011110000111100001111000011101100111011001110111011101110111011101111000011110000111100001111000011101100111011101111000011110000111100001111000011110000111011101110111011110000111100001111000011110000111100001111000011101100111011001111000011110000111011101110111011101100111011001110110011101100111100001111000011110000111100101111000011110000111100001111001011110110111110101111101011111011000001010011000100101101000111110011001101001111001000001010111101000101001010001011110010000100011001000100011011010110101101100110001001010110010101000100001,
	960'b000101110001111000100101001001100100011010000000001101000010110000111000010110011010110110111001010111111000100010100101100110001000111110011001100100010111111101111111011110110111110001111100011110000111100001111000011110000111100001111000011110000111011101111000011110000111011101111000011110000111100001111000011110010111100001111000011110000111011101111000011110000111011101110110011110000111100001111000011110000111100001110111011110000111011101110110011101110111100001111000011110000111100001110110011101110111100001110111011110000111100001110111011101110111100001111000011110000111011101110111011110000111011101111000011101110111011101110111011110000111100001111000011101100111011001110110011110000111100001111000011110000111100001111000011110000111100001111000011110110111110001111101011111010111111110000100100110111001010110010001100111001010100001111100011011001010010001111010010001010010111100100001001111110111010000111110001010010010011000100011,
	960'b000111000001111000100000001011100110000101101011001001000010101100111000100000111011110010001000011011111010010110011010100011111001100110010110100000000111111110000000011111010111101101111001011110000111100001111000011101110111011101111000011110010111100001110111011110000111100001111000011110000111100001111000011110000111100001111000011101110111011101110111011101100111100001111000011110010111100001111000011101110111011101110110011101110111011101110111011101100111011101111000011101110111011001110110011101110111100001110111011110000111100001111000011101110111100001111000011101110111011101111000011110000111011101110111011101110111011001110110011101110111011101110111011101100111011001110111011101100111011101111000011110000111100001111000011110000111100101111000011110000111100101111011011111000111111110000001100001111001111010010010100101001001111010100101011001011000111010010001010110000011001000100111000111100111000001010001001100010010011000100010,
	960'b000111010001111000100010001101110111011101000010001001010010100101001010101001001011001101100101100110001001110010010000100100001001101110000011011111110111111101111100011110100111100101110111011110000111100001111000011110000111100001111000011101100111010101111000011110000111100001111000011110000111100001110111011101110111100001111000011101110111011101110111011101100111100001111001011101100111011101110111011110000111011101110110011101110111011101110110011101100111100001111000011101100111011101110111011101110111100001111000011110000111100001111000011101110111100001110111011110000111100001111000011101110111100001111000011110000111100101110111011101110111011001110111011110000111011101110111011101110111011101111000011101110111100001111000011110000111011101111001011110000111100001111010011110110111111010000001100000101000110010011100100011101001010110100001100011110110100110011010011100110011101000100111000110100101000001100111001100100010011000100010,
	960'b000101110001111000100101010001010111101000100111001001100010101001101100101100001000110101110110100111111001010010001010100110101000101110000000011111010111110101111011011110010111100001111000011110000111100001111000011110000111100101111001011110000111011101110111011101110111100001111000011101110111011101110111011101110111100001110111011101110111011101111000011110000111011001110110011101100111011101110111011101110111011001110110011101100111010101110110011101100111011001110110011101010111011001110110011101100111011001110111011101100111011101110111011101100111011001110110011101110111011101111000011101110111011001110111011110000111011101110111011101100111011101111000011101110111100001110111011101110111011101110111011101110111100001111000011110010111100001111000011101110111100001111001011110110111110001111110100000001000000010010110100100111000101010010110101000000110111010001110100001110100101100101000001000000011000101101111001110100010100100100100,
	960'b000110000001111100100111010111000110010000011111001001000011010110001010101010110111000010010010100110001000110010001110100101101000000101111111011111010111101001111011011110100111100001111001011110000111100101111000011110000111011101110111011110000111100001111000011110000111011101110111011110010111100001110110011101110111100001111000011110000111100101110111011110000111011001110101011101110111011101110110011101010111011001110110011101010111010101110110011101010111011001110101011101100111010101110110011101100111011001110110011101000111011001110101011101100111010101110101011101110111011101110110011101110111011001110111011110000111011101110110011101100111100001111000011110000111100001110111011101110111011001110111011110000111011101111000011110000111100001111000011110000111100001111001011110110111101101111101011111110111111110000101100110111000100110001110100110101000101001110111100100100101111100101100001000110001101101101010010011010010100100100011,
	960'b000110010001110100101101011100000100011000011111001000100100100010011010100111010111001110011011100011011000010110010111100010010111110101111100011110110111101101111011011110100111100001111001011101110111011101111000011110000111011001110111011101110111011101110111011101110111011001110111011110000111011101110110011101100111011101110111011110000111011101110101011101010111010101110110011101100111011001110101011101100111010101110110011101100111011001110101011101010111011001110110011101100111010101110110011101100111010101110110011101100111010101110101011101100111011001110101011101100111011001110110011101100111011001110110011101100111011101110111011101110111011101111000011110000111011101110110011101110111100001110111011101100111011101111000011110000111100001111000011110000111100001111001011110110111101001111011011111000111110101111101100100101000111010000111100100001001011101110010100100000111001100110101001000100001011001010110010110100010101100100101,
	960'b000101110001110100110111011101000010101100100000001001100101110010011110100010011000011010010101100010001000100010010100011111000111100101111010011110110111101001111011011110100111100001111000011110010111011101111000011110000111100001111000011101110111011001110111011101110111011101110111011110000111100001110111011101110111011001110110011101100111011001110101011101010111010101110110011101010111011001110110011101010111011001110110011101100111010101110110011101100111010101110101011101100111011001110110011101010111011001110110011101100111010101110101011101010111011001110110011101100111010101110101011101100111010101110110011101010111011001111000011110000111100001110111011101110111100001110111011101100111100001111000011101100111011001111000011110000111100001111000011110000111011101111000011110010111101001111010011110110111110001111100100001101001001110000011100010011001011001111101100010011000000001000010001000110001100000111001011001000011001100100100,
	960'b000110000010000101000101011011010001111000100010001010110110110110011100011111111000111110001100100001001000110010001010011110110111101001111011011110110111011101111000011110010111100101111001011110010111100101111000011110000111011101110111011101110111011101110111011101110111011001110111011110000111011101110111011101110111011001110110011101100111011001110111011101110111011001110101011101010111011001110101011101100111011001110110011101100111011001110110011101010111011001110101011101100111010101110101011101100111011001110110011101010111011001110110011101100111010101110110011101010111011001110101011101100111010101110110011101100111011001110110011110000111100001111000011110000111011101110111011101100111100001110111011110000111011101110111011110000111100001111000011110010111100101111001011110010111101001111001011110010111101001111011011111101001010110000011100001101001000010001100100000001000011101001111001001100001110000100110011001110011100100100100,
	960'b000110010001111101001011010111100001101000100010001100100111011110010101100000001001001110001010100000011001000010000100011111000111101001111010011110010111011101111001011110000111100001111000011110000111100001111001011101110111011101111000011110000111100001110110011101100111011101110110011110000111011101110111011110000111011001110101011101010111011001110111011101110111011001110101011101100111011001110110011101100111011001110110011101100111011001110101011101110111011101110110011101100111011001110101011101010111010001110101011101010111011101110111011101100111010101110110011101010111011001110110011101100111010101110110011101000111011001110110011110010111100101111000011110000111100101110111011101110111100001110111011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111001011110010111100101111010011111001000111110000111100001001000101110010010100000011000100101011100001010100010000100011011011000010011110000100100,
	960'b000110100010001001010011010011000001110000100101001110110111101110010001100001111001010010001000100000001001001010000000011110110111101001111000011101110111100101111000011110000111011001110111011110000111100001111001011101110111100001110111011110000111100001110111011101100111011101110111011110000111100001110111011110000111010101110101011101100111011001110110011101010111010101110110011101010111010101110110011101100111010101110110011101100111010101110110011101100111011101110110011101100111011001110110011101010111011001110111011101100111011001110101011101100111010101110110011101010111010101110101011101100111011101110111011101100111011001110111011110000111100001111000011110000111011101110111011101110111011101110111011101110111100001111000011110000111100001111000011110000111100001111001011110000111100101111000011110100111100101111010011110111000100010001100100000001000100110010100100001101000101101100100001011100010001100011000010110000100010000100010,
	960'b000101100010010101011001001111000001111000100111010000010111110110001101100011101001010010000111100000011001010001111110011110100111100101111010011110100111100101111010011110000111100101111000011110010111100001111001011110000111100101111000011110000111100001111001011101110111011101111000011110000111100101110111011101110111011001110110011101010111011001110110011101010111010101110110011101100111010101110110011101110111010101110101011101010111010101110101011101010111011001110101011101100111011101110101011101100111011001111000011101100111011001110110011101010111010101110101011101010111011001110110011101100111100001111000011101010111011001110110011101110111011101110110011101100111011001110110011101100111011101110111011101110111100001110111011101110111100001111000011110000111011101111000011110010111100001111000011110100111101001111010011110111000010110010000011111111000100010010111100011011000110001101010001101010010010000010110010011100100100100100011,
	960'b000110000010001001011001001100100001111100101010010001100111101110001011100101101001010010000111100001011001001101111100011110110111101101111011011110100111100101111001011110000111100001111000011110000111100001111000011110000111100001111000011110000111011101111001011101110111100001111000011101110111100001111001011101110111011101110101011101000111010101110111011101010111010101110110011101010111011001110101011101100111010101110110011101100111010101110101011101100111011001110101011101010111011001110101011101100111100001110110011101100111100001110110011101100111011001110110011101100111011001110111011110000111010101110110011101110111010101110101011101110111011101110110011101110111011101110110011101110111100101111001011101110111011101110111011110000111011101111000011110000111100001111000011110000111100001111000011110110111101001111101011110101000001110010010100000101000100110010110100101011000110001101100001110010010011100011000010001100100110000100010,
	960'b000110110010011101011001001011110010000100101101010001110111100110001111100111001001011010001001100001111001001101111101011111010111110001111010011110110111101001111001011110000111100101111000011101110111100001111000011101110111011101111001011110000111100001111000011101110111011001110111011101100111011101110110011101100111010101110110011101010111011001110101011101100111011001110101011101100111011001110111011101110111010101110110011101010111011001110101011101010111011001110101011101010111010101110110011101100111010101110101011101100111011001110101011101010111011001110110011101100111010101110101011101010111011001110100011101010111011001110111011101100111011101110110011101110111011001110110011101100111011101111000011101110111100001111000011101110111100001111000011110000111100101110111011110000111100101111001011110100111101001111100011111101000001110010101100001001000101110011000100111001000110101101101001111000010100100011000010010000100110100100100,
	960'b000110010010010001011011001100010010001000110000010010000111011010010011101001001001100110001101100010101001011001111111011111100111101101111011011110010111101001111000011110000111100001111000011110000111100101111000011110000111011001111000011110000111100001110111011101110111011101110111011101100111011101110111011110000111011101110110011101010111011001110110011101010111010101110110011101100111011001110111011101100111010101110110011101100111011001110110011101100111010101110101011101100111011001110110011101100111010101110110011101100111010101110101011101100111010101110101011101100111011001110101011101010111011001110101011101010111011001110111011101110111011101110110011101100111011101110110011101110111100001111000011101110111100001111000011101110111100101111000011110000111100001111000011110010111100001111010011110110111110001111101011111111000010010010110100001111000111010011100101001011001000001101100001111110010101100011011010001110100110100100110,
	960'b000101110010011001011011001100100010001100110011010010100111001010001111101010101001111010010001100011011001100010000100100000000111111001111101011110010111100101111001011101110111100001111001011110010111100001111000011110000111011101110111011110000111011001111000011110000111011101110111011101110111011101111001011110010111011101110111011101110111011001110111011101100111010101110110011101110111011101110110011101010111010101110110011101100111010101110111011101110111011001110111011101100111011001110110011101010111011101110111011110000111010101110101011101010111011001110111011101010111010101110101011101000111011101110111011101110111011101110111011101100111011101111000011110000111100001110111011101110111100001110111011101110111100001111000011110000111100101110111011110000111100001111000011110010111100101111010011110110111110110000000100000011000101010010111100010111001010010100000101010011000111001101010010000010010111100011100010010000100111100100010,
	960'b000110000010010001010111001101000010011000110111010011010110110110001011101011101010010110010111100100001001101010000111100000010111111101111101011110110111101101111011011110000111100001110111011110000111100001111000011110000111100001111000011101110111011101111001011101110111011101111000011101110111011101110111011101100111011101111000011110010111011101111000011110000111011101110101011101100111011101110101011101010111011001110110011101010111011001111000011101110111011101110111011110000111100001110110011101110111011101110111011101100111011101110110011101100111011001110110011101010111011001110110011101110111011001110111011110000111100001110111011101110111100001111000011110000111100001110111011101100111100001111000011110000111011101111000011110010111100001111000011110010111100101111000011110000111110001111010011110110111110110000000100000101000111110011010100011111001100110101000101011111000101001100100010001000011000100011100010010100100101100100111,
	960'b000110000010010001010110001101100010100100111100010100110110011110000101101100111010110010011100100100111001111010001100100001001000001001111111011111010111101101111010011110010111100001111000011110000111100001111001011110000111100001111000011101110111100001111001011101110111011101110111011110000111011101111000011101110111011101110111011110000111100001110111011101110111100001111000011101110111011101111000011110000111011101111000011101110111100001110111011101110111011101110111011101100111011101111000011101110111100001110111011101110111100001110111011101110111100001111000011101110111011101110111011110000111011101110111011101110111011101111000011101110111011101111000011110000111011101110111011101110111011101111000011101110111100001111001011110000111011101111000011110000111100001111001011110010111101101111101011111101000000010000011100001001001100010011001100101001001111110110000101100001000010001100000010011000011011000011110010011000100110000100110,
	960'b000101100010010001010111001110110010110001000011010110110110000001111110101011111011010010100100100101111001111010010100100001011000010010000000011111010111101101111011011110110111100101111001011110000111100001111001011110000111100001111000011110000111100001110111011110000111011101110110011110000111100001111000011101110111011001110111011110000111100001110110011101110111100001111000011110000111100001111000011110000111100101111000011101110111100001111000011110010111100001111001011110000111100001111000011110000111100001111001011110000111100001111000011110000111100001111000011110000111100001111000011101110111100001111000011110000111011101111000011110000111100001111000011101110111100001111000011110000111011101111000011101110111100001111000011101110111100001111000011110010111100001111001011110010111101001111110011111111000001010000110100010011001111010011000100110111010011110111001101010110111110001011100010101100011100100100011010011010100111000100110,
	960'b000101100010000101010011001111110011001001001001011001100101110101110101101000111011111010101010100111001001110010011101100010001000010010000000011111110111110001111011011110010111100001111001011110000111100001111000011110000111100001111000011110000111100001110111011110000111011101110111011110000111100001110111011101110111100001110111011110000111100001111000011101110111100001111000011110000111100101111000011110010111100001111000011110010111100101111001011110010111100101111010011110010111100001111000011110010111100101111001011110100111100101111001011110010111100101111001011110000111100001111000011110000111100001111001011110000111100001111000011110000111100001111000011110000111100001110111011110000111100001111000011101110111100001111001011110000111100001111000011110000111100001111001011110100111101101111110100000011000010010001000100011011010001110011001101000011010111010111111100111010111010001100000011000010011111000101000010100010100011000100011,
	960'b000110010010000001001100010001100011100101010000011100000110010101101101100100011100001010110001101001001001100110100011100011001000011010000010011111110111110101111011011110010111100001111001011110000111011101111000011110000111100001111000011110010111011101111000011110000111011101110110011110000111100001111000011110000111011101111000011110000111100101111001011110010111100101111000011110000111100101111001011110010111100001111001011110010111100101111011011110110111101001111010011110110111100101111010011110110111101001111010011110100111101101111001011110000111101001111010011110000111100101111001011110010111100001111000011110000111100001111000011101110111100001110111011101110111100101111000011101110111011101111000011101110111100001111000011110000111100001111000011110000111100101111011011110110111101101111111100000011000011010001000100110001010001010011001101001011011011011000001100011010110100101110001011010010100001100101101010101100011111000100011,
	960'b000110010001111101000101010010010011111001011000011101000111100101100100011111111011100110111001101010001001100110100001100101111000011010000100100000000111110001111011011110110111100001111001011110000111100001111000011110000111100001111000011110000111100001111000011110000111011101110111011101110111100001111000011110000111011101111000011110010111100001111000011110010111100101111000011110010111101001111001011110100111101001111010011110100111101001111100011110110111101101111011011111000111110001111100011110110111110001111100011110110111101101111010011110100111101101111010011110100111100101111010011110010111100001111001011110010111100001111000011110010111100001111000011101110111011101111000011101110111011101111000011110000111100001111000011110000111100001111000011110000111100101111010011110110111110101111111100000101000011110001011101000111001101110011110101010111011111010110100011111010110001110000100011011000100100000110010010110100011101000011100,
	960'b000101110001111101000001010100010011111001011101011101001000101001011111011101011010010011000001101011011001111010011000101000011000100110000100100000010111110101111011011110110111100101111001011110010111100001111000011110000111100001111000011110000111011101111000011110000111100001111000011101110111011001111000011110000111100001111000011110000111100001111000011110000111100101111000011110010111101001111010011110110111101101111011011111000111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111100011111000111110001111011011110110111101001111011011110110111100101111001011110100111100101111001011110000111100001111000011110000111011101111000011110000111100001111001011110000111100001111000011101110111100001111000011110000111100101111010011110110111110001111111100001001000011110010100101000101001100010100100101100011100010010011001011100010110110110001100011010100100110100110011010110100011010000100010,
	960'b000110110001110100110100010110010011001001100000011100101000111101101101011010111000100110111101101101001010001010010110100110111001010010000010100000010111110101111011011110100111100001111001011110010111100101111000011110000111100001111001011110000111100001111001011110000111100001111000011110000111011101110111011110000111100001111000011110100111101001111001011110010111101001111011011110100111101101111100011111000111110001111100011111100111111101111110011111111000000010000000100000000111111110000000100000001000000010000000011111110111111001111110011111100111110101111100011111000111110001111100011110110111101101111011011110100111100101111000011110000111100001111000011110010111101001111001011110010111100001111000011110000111100101111001011110000111100001111001011110010111100001111010011110110111110001111110100000111000011110011111100110001001110010100111101110011011100110000000011000101000100110001001011001100100111100110101010111000010110100100001,
	960'b000111000001111000101011010111010010110001011011011011001000010110001001010111000111011110100110101110111010010110011000100011111001110110001001011111110111111001111011011110100111100101111001011110010111100101111001011110000111100101111001011110010111100101111000011110010111100101111010011110010111100001111001011110010111100101111001011110010111100101111010011110110111101101111011011111010111110101111110011111110111111101111111011111101000000010000001100000001000000110000010100000011000001010000010100000111000000110000001100000011000000110000001100000010111111101111111011111110111111101111110011111010111110001111100011110110111101101111010011110100111100101111001011110100111101001111010011110100111100001111010011110100111101001111010011110100111100101111001011110010111101001111010011110110111110001111111100000101001010010011010100100111001111010101101101111111001101001110010011001101001001101111000010110110100000001000010010100110010100000100001,
	960'b000110000001111000101001010100110011101101000001011001100111001110010010011010000110101110000101101101111010110110011100100100001001000010011001100000010111110001111101011110110111100101111001011110100111101101111010011110100111101001111010011110110111101001111010011110100111101001111010011110010111101001111001011110010111101101111100011110110111101101111100011111000111110001111101100000001000000010000001100000011000000010000000100000101000010010000100100001001000010010000100100001011000010110000101100001001000010110000100100001001000001110000100100001001000000110000001100000011000000110000001100000000111111001111101011111010111110001111100011110110111110001111100011110110111101001111011011110110111100101111010011110100111101101111011011111000111101001111010011110100111101101111011011110110111111010000001100011101001100110001100100101101001111110110011101100100111111001100011011110010111111001100101010110000010100001010101010001000010101000100011,
	960'b000110010010000000100101010001000101010100011111010111010110000001111111100001100101100001110111100110001011000110100000100100101000100010001101100101000111111101111100011110110111101001111011011111000111101001111011011111010111110101111110011111010111110001111101011111010111101101111011011111000111110101111010011110100111101101111101011111100111111001111101011111110111111110000000100000001000001010000010100000111000010010000100100001011000011010000110100001111000011110000110100001101000100010001001100001111000011110001000100001101000011110000110100001011000010110000101100001001000010010000100100000101000000110000000011111100111111001111111011111010111110001111100011111000111110101111100011111000111101101111100011111010111110101111101011111010111110001111100011110110111101101111011011111100111110110001000100110001000100110001101100110001010010110110101100011110111000001011011011110000110001101010001010010100010000101100010001110100010011100100011,
	960'b000110100001111000100100001110110110000100100000010000000101000001011110011110010110001101100100011111011010001010100110100110001000110110000100100011001001010010000000011110110111110001111100011111000111110001111101011111110111111101111111011111110111111101111110011111100111111001111110011111010111110101111011011111000111110001111101011111101000000010000000100000011000001110000100100000111000010110000101100001111000010110000111100010001000100110001001100010101000100110001010100010101000101010001010100010111000101010001010100010011000101010001000100010001000100010001000100001011000010010000100100001001000001110000010100000011000000001111110011111110111111001111101011111010111110101111101011111100111111101111111011111110111111101111111100000000111111110000000011111100111110101111110011111101000100110010101100001111000100010001111100111011010101010011001011101110101101101011111010110110100101101001101001001100011110101011100001100000010010100100111,
	960'b000110000001111100100101001100100101011001000100000101110100100101000110010101010110110001010010011011101000010110100110100111111001001110001010100000111000100110010101100001100111110001111101011111010111111110000000100000001000000110000001100000111000001110000011100000101000000110000000011111110111111101111110011111100111111001111111011111100111111110000011100000111000010010000110100001011000011010000111100010001000100110001010100010101000101010001100100011001000110110001101100011011000110110001110100011011000110110001110100011011000110110001011100010111000101010001000100010101000100110000111100001111000010110000100100001001000001010000001100000000111111101111110011111100111111010000000100000001000001010000010100000111000001010000011100000111000000110000010100000001000000010000010100011111001010110000011100001001000110110011001101001011001110001111011011001110100111101001111010000000011101100111110000100010101110101000111001010110010101000100110,
	960'b000110000010000100101000001010110100011001100011000101010010111101000011010000010100111001010111010011110111001110001010101001001001110110010010100010011000001010000100100100101001001110000111100000011000001010000011100001001000010110000101100001101000011010000101100001001000010010000011100000011000000110000010100000011000000110000010100000101000001010000011100001011000010010000111100010001000100010001010100010111000110110001100100011101000111110001111100100001001001010010000100100011001000110010001100100011001001010010001100011101000111010001110100011011000110110001100100010111000101010001001100010011000011110000111100001111000010110000011100000111000001110000010100001001000001010000011100001001000010110000101100001101000011010000110100001011000010010000100100001101000111110010111100100001000010010000111100011011001010010100000101000010111111101101110010010000100001100110110001100000011110000011001001011010110001100110111001010110010110100100101,
	960'b000110010001111000100101001011100011001001011100001111100000110000111011001101100011110101000111010011000101001101110101100011011010001010011011100100101000101110000110100000111000110010010111100101111001001010001101100010101000100010001000100010101000101010001001100001111000100010000110100001101000010010000011100001001000010110000100100001001000010110000110100001111000100010001010100010111000110010001110100011101001000010010000100100011001000110010010100100101001001010010010100100111001001110010010100100101001010010010011100100011001000110010000100100001000111110010000100011101000111010001011100010111000101010001010100010101000011110000110100001001000010110000100100000111000011010000110100001111000100010001001100010101000101010001010100011001001000110011000100111011001100110001011100010001000101110001111100101111010000110100000100000000111000101001010001111010010111000101011001011110010100100001101010110100100110000110011001011010010011100100101,
	960'b000110010001111100100100001011000010101101000101011001010001011000011010001110000011000100111000010000010100011001010100011101101000110010100011100111101001011110010000100011011000101110001011100100001001100010011111101000001010000010011111101000001010000110100000100111101010000010011011100110101001100110011000100110001001100110011000100110011001101010011011100110111001111010011111100111111010000010100001101000101010001010100011101001001010010010100101101001011010010110100110101001101010011010100110101001101010010010100101101001011010010110100100101001001010010010100010101000101010000110100000101000001001111110011100100111011001110010011011100110011001100110011010100110001001101110011011100111001001110110011110100111111010000010100001101000111010001010011100100101011000111110010001100100101001011110011011101001001001110001111111011100010100011100110011001010110010100000100011001011000000110000110110011000110011101100110000001011100010011100100100,
	960'b000101110001111100100100001010000010111100111010010110110100011100001001001001000011001100110000001110000011100100111111010011100111000010000111101000111010010010011011100110011001011110010110100101011001011010011000100110111001111010011101100111101001110110011011100110111001101010011000100101011001001110010001100100101001000110010001100100111001010110010100100101101001100010011001100110111001110110011100100111011001111010100001101000001010001010100001101000101010001010100010101000101010001110100010101000101010000110100010101000101010000010100000101000011001111110011101100111101001110010011011100110011001101010011001100101101001010110010101100101001001010010010100100101001001010010010111100110001001100110011100100111001001110110011110100111011001110010011100100111011001110110011110101000011010010110100110100101000111110001101101010000110010110000101001001010000010000100101000000100100001011001011111010100100011110000101111001011010010101000100100,
	960'b000110010001110000100100001001110011000100110001010000110110100000101001000010010010100100101111001011110011001100110100001111010100100101100111011111101001101110101011101010011010001110100010101000111010010010100110101001101010011010100111101001111010011110100101101001011010001110100000100111101001101110011001100110001001100010011000100110011001101110011011100111101001111110100000101000101010010010100011101001101010010110100111101010001010011110101000101010011010100010101000101010001010100110101000101010001010100110101001101010001010100010100111101001111010011110101000101001101010010010100011101000111010000010100000100111011001110110011010100110101001100110011001100111001001110110011111101000001010010010100101101001101010100010101001101010111010101110101010101011011010111010110001101100001010001110001001011101110110001000111101001010100010010100100101000111100010011000010110000011000100101101100011001111110011011000110011001010100010011000100011,
	960'b000110110010000000100011001010010010101100110011001111000101010101100010000101000000110000101100001011110010111000110011001101010100000101001000010110010111000010000111101001011011011110111001101101111011100010110111101101111011011110111000101101111011011110110110101101001011001110110000101011101010101110101000101001111010011110100110101001101010100010101001101011001010110010101110101100001011000110110010101100111011010010110100101101001011010110110110101101101011011110110111101101101011011110110110101101101011011110110110101101001011010110110100101101011011001110110100101100111011001010110000101100001010111010101101101011001010101010101001101001111010100010101001101010101010101110101110101100001011001010110101101101111011100010111010101111001011111010111111110000011011110010101011100100010111110101101101010100000011011000101010001001110010001000011100001001010001100100001010001100010110110101001100001101110011011000110100001011110010100000100011,
	960'b000110100001111000100101001010000010110100110000001101110100000101100010010100110000110000001110001011000011001000101011001011110011000100111111010011110101000001011101011011101000001010011100101100101011111111000110110010111100110011001110110011101100110111001100110010011100100011000101110000111100000110111110101111011011110010111100101111011011110110111111110000001100000111000011110001001100010111000110110001101100011111000111110001111100100011001000110010001100100011001000110001111100100111001001110010001100100111001000110010001100100111001000110010011100011111000110110001101100011011000101110001001100001011000011110000101011111011000000101111111011110110111101101111111100001011000011110001011100011111001001110010111100110011001011110010101100011010110110101000111000110001111011011010110101011101000011001101100010100100100101001000010001111100101000000110100000101100100001011010000100111000111011001110100011100000110011001010110010100000100011,
	960'b000101110001111100100101001010000011000000110100001100010011101101001000011001000100010000001100000011010010011100110111001001110010101100110000001110000100100101010110010101010101011101100001011011110111110010001011100101101001111010100011101001101010100010101001101010101010110110101111101100001011000110110010101101001011010110110110101101111011100010111010101110111011101110111101101111101011111010111111110000001100000011000001110000011100000111000010110000101100001011000010110000111100001111000010110000111100001111000011110001001100010011000011110000101100001011000010110000101100000111000001101111111011110110111011101110101011011110110110101101001011000110110000101011011010101010101000101001111010010110100011101000101001111110011000100100001000010001111001011011100110000101010010010001100100000000110100001010000010001100100000001000110010110000010111000011000001100001011110010110110100000000110011001110010011100000101111001011100010101000100010,
	960'b000110100001111100100100001011010010110100110011001101110011010000111001010001000110110001000000000010110000110000011100001101110010110000100110001011000010111000110111010001010100111001010001010100110101011101011010010111100110000001100010011000110110010101100110011010000110100101101001011010100110110001101101011011100110111101110000011100100111001101110100011101010111010101110111011110000111100101111011011110100111101101111100011111010111111001111110011111101000000010000000100000001000000001111111011111111000000001111111100000011000000001111111011111100111111001111100011110110111101001111000011101110111011001110101011101000111000101101111011011100110110001101010011010100110011101100110011001100110010001100011011000110110001001100001010111100101100001010000010010010100010001000000001100110010101100100111001001000010000100101011001010100001001000001110000101100101101001100100001111000011100000111001001100100011000100110001001011010010010100100101,
	960'b000110100001110100100100001011100010110100101111001101110011011000110110001111000100100101101000010000010000111000001011000100110010111000110011001010000010010100101011001011000010111000110101010000000100101001001011010010010100101001001001010010010100100001000110010001100100001100111111001111010011110000111100001111010011110100111101001111110100001001000011010001010100100001001010010011100101000001010001010100100101011001011000010111100101111101100000011000000110000001100000011000000110000101011101010111010101101001011011010111000101101001011000010101100101010001001111010010110100100101000110010000110100001101000001010000110100001101000011010000110100001101000011010001110100011101001000010010100100101001001001010010010100101101001100010010110100011000111100001101010010111000101001001001100010010100100100001010010010111100100000000011100000110100011010010110010110000101000100001101100011010000111001001100110011000100110011001010110010011100100101,
	960'b000110000010000000100110001010010011000100110010001100110011010000110101001101100011100001001101011010110100101100010011000011000000110100011010001100100011011100101101001000110010001100101000001010100010111000101101001011110011000000101110001011110010111100101110001011010010101100101001001010010010100000101000001010000010011100100110001001110010011100101001001010110010110000101010001011000010111000110000001100100011001100110100001101010011011000110110001110000011100100111010001110110011110000111011001110110011101000111001001101110011010100110101001100110011000100101110001011000010110100101100001010010010100100101000001001110010011100100111001001110010011100100111001001110010101000101101001011110011000100110010001100110011001000101111001100000010110100101010001010100010100000100110001010000011000000110100001001110001001000001101000011000010000001011111011001100100010000111001010000000011101000110010001100110011001100101110001010110010110100100101,
	960'b000110000010000000100101001010110010111100110010001100110011010000110011001110000011011100111011010001100110011001011011001000010000110000001101000011100001111000111001010000110011101100101100001000110010001000100011001001100010011100101001001010010010101000101010001010000010100000100111001001110010011100100110001001010010001100100011001000100010000100100011001001010010011000100110001001100010100000101011001010100010101000101010001010100010110000101101001011100010111100101111001100000011000000101111001100000011000000101110001011000010101100101100001010100010100000100110001001110010100000101000001010000010011100100111001001100010011000100110001001010010010000100100001000110010010100100110001001010010010100100101001001110010100000101000001001110010010100100101001011000011011101000001001111100010101100010011000010110000101100001110001100110110011101011000001111110011101000111010001101110011011000110110001100100011000100110010001010110010100000100100,
	960'b000110100001110100100101001011110010101100101110001101100011010100110101001101110011100100110011001110110100100101011010011001110011111000010011000011000000110000001111001000010100011001100010011000110101011101001111010011100100111001001111010011110100111101001110010011000100101001001011010010110100101001000110010001010100010001000100010001010100010001000011010001010100011001000110010001110100011101001000010001110100100101001001010010110100101101001101010011110101000001010000010100010101001001010001010100010101000001001111010011000100101101001001010001110100011101000101010001000100010001000010010000010100001001000010001111110100000001000010010000110100010001000011010001000100001101000100010001010100010101000100010001110100011101000101010001100100111101011000010101110100001100100111000101000000110000001110000100000001111001001111011010100101000000111101001100100011011000111100001100100011010100111010001100100011000100110000001011010010010100100101,
	960'b000110100010000000100100001010010010101100110011001101000011010100111010001100110011101000111000001101100011100100111010010100000110011001011101001100010001000100001100000010110000110000011001001100000100010001001000010001110100101001001001010010110100110001001010010010110100100001001000010010000100011101000111010001100100010101000110010000100100010001000100010001010100011001000111010010000100100001001010010010000100101101001110010100000101001001010100010101110101100001011000010101110101101001011011010110010101100001010110010100110101000001001101010010100100100001000111010001100100011001000011010000100100000101000001010000100100000101000100010001010100011001001000010010010100101101001010010010110100110001001011010010110100110001001001010010010100000100101101000110000000111000001101000011110001000100011101010001000110011001011111010001110011100000110111001110010011001100110101001101100011100100110110001101100011010000101100001011110010100100100001,
	960'b000110000001111100100101001001100010110100110010001100000011101100111101001101100011010000111001001110000011010000111001001110000011111001011101011011010101110100111000000111010000111100001100000011000000110000001010001011001010100101011101000010100000110100010000100001001001000100010111000011110000111100001111000011010001100010010100100000100001000100001110000011100000110100001110000011010001011110010100100000100001000100001110000011110000111100001101000011010000111110000010100100010001011100001101000011100000111000001110000011100000110001110010100111110010000100001101000011100000111000001110000011100000101001011111101010000010110100001010000011010000110100001101000011111000001110010001000101100000110000001000010010111010101100111000000010010000110100001100000011010001000000010101001010000100011101100101011000100100101001000000001110110011101100110101001101110011100100110011001110010011011100110100001110110011100100110000001010010010100000100011,
	960'b000110100001110100100010001001110010101100101111001101110011011100111001001110100011100100110100001101100011011100110100001101100011110100111101010001110101100001101001011001010101000000111001001001100001101000010011000111110110110101000101000011110001000100010010010100100110011000010110000100000001000000010001000100000001010001011011010111010001000100001111000011110000111100001111000011110001001101011011010110110000111100001110000011100000110100001101000010110000111001010000011001100001000100001011000010110000110000001100000011000000110101000100011011100001101000001101000011000000110100001110000011110000111000111001011100100010001000001101000100000000111100010000000100100101000001100111000101100001000100010001001011110111001100101111000100100001100000100000001011100100011101011110011010000110000101001011001111110011110000111001001110100011101100111011001101100011010000110101001101100011100000111100001101110011011000110011001011010010011000100010,
	960'b000111000001111000100001001010000010100100110001001110010011011000111001001110110011110000110110001101100011011100110111001110100011111100110111001110010011110101000011010010010101100001100100011010010110010101011111010101000100110101001101010011010100111101001111010010110100100101001110010011100100111101001110010011110100110101001010010010110100111001001100010100000100111001001111010011100100110101001000010001110100110101001100010011010100111101001110010011010100111001001001010001100100101101001110010011010100110001001110010011010100110001001100010010000100110001001110010011000100101101001101010011010100110001001011010010100100110001001110010011100100110101001101010100000100101101001010010011100100110101001111010011100100101001001111010110000110001001100111011010100110010101010010010001000011110000111000001101010011110100111001001110010011101000111100001101100011010100110110001101110011011100111100001101110011010100110010001011000010011000100011,
	960'b000101110001110000100011001001100010100100101110001100100011101100111010001110000011010100111000001110000011100000111010001101100011011100111110001111000011100100110011001110000011110000111101010000110100100101010100010110110101111001011100010110110101110001011011010111000101110101011010010111100110000101100000010110100101110001011101010111010110000001011100010110100110000101100000010111010101100101011010010111010101110101011110010110110101110001100010011000010101111001011001010111000101110001011100010111000101101101011011011000110110000101011011010110100101111001011101010111100101110001011000010111000110000101100000010110100101110001011001010101110101101101011011010111000110001001100000010110100101111001011101010111000101110101011011010101000101001101001111010001100011100100111010001110100011011000111001001101110011001100111100001110110011101000110100001110010011011100110110001110010011011100110011001111000011100000101111001011000010100100100100,
	960'b000110000001111100100001001001010010100100110010001100100011010100111100001101100011100100111010001101100011100000111001001110100011011100111011001111000011010000111001001110100011100000110101001110010011100000110101001111000011101100111000001111010011101100111000001110010011110000111011001110100100000000111001001110010011110100111001001110010011101100111101001110100011110000111111001101110011101000111100001110000011100000111100001110110011011000111110001111100011100000111010001111000011011100111000001110010011101000111000001111100011101100111000001110110011101000110110001101100011100100111001001110000011111000111000001110000011011100110110001101010011011100111010001110000011101000111010001110110011110100111000001110100011100100111011001110110011011100111101001101000011011100111010001101110011100100110111001110100011011000110110001110010011011000111001001110010011011000111000001101110011100100110110001101010011010100101111001011110010100000100011,
	960'b000110010001110000100011001011000010101000101110001101010011010000110110001101100011101100110110001110100011111000110111001101110011101000110110001110010011011100111001001101010011110000111100001101010011100100111000001101110011010000111001001110000011010100111110001110100011011000111001001101110011100000110100001110100011011000111001001111100011011100110110001110100011010100111001001101010011101000110110001110010011101100110101001101110011100000110101001101100011010100111001001101010011100100111011001101000011010100111000001101010011010100110111001101110011010000111011001110100011001000110111001101010011011000110011001110010011001100111000001110000011000100110111001101110011011000110110001110100011011000110101001111000011101000110101001110100011100000111000001101100011101000110110001110000011111100111000001101100011101100110111001101110011011000111011001101010011100000111101001101110011011100111010001101000011001000110001001011010010011000100111,
	960'b000110000001110000100010001010100010101100101111001101000011010000110100001110100011011100111001001110010011101100110111001101100011101000110100001101000011100000110101001101010011101100111011001101110011011000111000001101000011010000111001001101010011011000111011001110010011011100110110001110000011010000110111001110010011011000111000001111010011100100110110001101110011011000110011001110000011011100110110001110000011110100110111001101010011011000110011001100100011100000110111001101110011100100111010001110000011011000111000001101000011010100111000001101100011100000111000001110000011011000110100001101010011000000110011001101110011011000110110001101100011100000110111001101110011010100110110001110010011100000111010001110000011100100111001001110000011011100110010001101010011011000110111001110000011101100111001001110010011011000110110001101010011011000110110001110000011100000111010001110010011011100110111001101000011000100110001001010110010101100100101,
	960'b000101110010000100100110001010000011000000110011001100000011001100111001001101010011010100111101001110110011100000111111001110110011011000110011001101100011010000110101001111000011100100111000001111110011011100110011001101110011100000110110001110100011111000111010001110110011110100110101001100110011100100110111001101100011110000111110001101110011111000111101001101000011010000111000001101010011010100111101001110010011011000111110001110010011010000110011001110000011011100110110001111010011101100111000001111010011100100110100001101010011011100110100001101110011111100110110001110010011111000110101001100110011011000110100001101000011101100110111001101110011101100110101001101000011100000110111001101100011100000111100001101110011101000111100001101100011010000110101001101010011010000111001001111000011011100111101001111010011010100110101001110000011011000110101001111110011110000111001001111010011100100110100001101000011001100101111001010110010110100100101,
	960'b000101110001110100100010001010100010110000101110001100100011010000110101001110000011011100110111001110000011101100111000001101100011100000110100001101000011100000110101001101110011101000111010001110010011011000111001001101000011011000111001001101010011011100111010001110000011100000110110001101110011010000111000001110010011011100111000001110110011011100110111001110000011011100110011001110000011011100110111001101110011101000110111001101010011100000110101001101100011100000110111001101110011011100111011001101100011010000111001001101010011010000111000001101010011011000111011001101100011010000110100001101100011001000110100001110000011010000110111001110000011010000110011001101110011010100110110001110100011011000110110001111010011100100110111001110000011011000110011001101100011100000110101001101110011111000110111001101100011100100110111001101100011100000111000001101100011011100111100001101110011011000110111001100110011001000110011001011000010011100100011,
	960'b000110010001110100100001001010110010100100101100001100100011000000110010001100110011100100110101001110000011101100110100001101110011011000110011001101000011010000110111001100010011100100111001001100110011100100110110001101010011010100111000001110000011010100111010001101110011001100110111001100110011011000110010001110100011010100110101001111000011010000110110001110010011010000110110001101000011100000110010001101100011100100110001001101010011010100110001001101010011010000111000001100100011010100111001001100100011011000110110001101000011001100110100001101100011001000111010001101010011000000110110001100100011010000101111001101010011001100110101001101100011001000110111001100110011001000110001001101110011011100110101001110100011010100110101001110000011000100110101001100000011011100110101001100110011101000110100001101100011100000110011001110010011010100111001001101010011010100111010001100110011011000110100001100010011000100101110001011010010011000100011,
	960'b000101110001111000100000001001010010100100101110001011010011001100110110001100100011010000110110001100110011001100110101001101010011001000110110001101010011000000110100001101000011001000110001001101010011010100110010001110010011100000110010001101100011010000110010001100010011011000110100001100110011100000110011001100100011011000110011001100100011001100110110001100100011011100111001001100110011010000110110001100010011000000110010001101010010111100111000001110010011001100110011001101010011000000110001001101000011011000110000001101100011011000101111001100110011001100101111001100000011010000110001001100010011011100110011001100010011010100110010001100100011010100110100001100110011100000110111001100000011010100110100001100010011001100110110001100100011010100110111001101000011000000110101001101010011000100110101001101100011000000111000001110100011011000110011001101100011010100110010001101000011010000101111001101100011010100101010001010100010011100100000,
	960'b000101100001101000100000001000110010100100101001001011000011001100110100001100110010111100110001001100000011000000110010001011110011000100110011001101000011000100101101001100010011000000110000001100100010111000110011001101100011011100110010001011100011000100110000001100010010111100101111001101000011010100110100001100000011000000110000001011110011001000101110001100010011010100110100001100110010111100110000001100010010111100110001001011010011000100110100001101010011010000101110001011110011000100110000001011110010111000110001001101000011010000110010001011100010111100101100001100000010111000101111001100100011001100110010001100000011000100101111001100000011000000110001001100110011010000110100001100110011000000110001001011110011000100101110001100100011001000110011001100110011001000101101001100010010111100110001001011110011001000110100001101000011010000110001001011110011000100110000001100000010111100110010001100010011000000101101001001100010001100011110,
	960'b000101110001101000011101001000100010010100101010001011110010110000101110001011110011001000101111001010110010110000101111001100100011001100101100001011100011000100110001001011010010110000101100001011010011001100110000001011100010111100110100001011110010110100101110001011000010111100110100001100010011000000101111001100110011000000101011001011010010101100110000001100010010111000101110001100010011010000101110001010100010101100101011001100010011000000101101001011100010111100110010001011010010110000101011001011000011000100110010001011010010110100110010001100100010110000101011001010010010110000110001001011110010110100101101001100000010111000101101001011000010111100110011001100000010111000101111001100010011000100101100001011000010110000101111001101000010111100101110001011110011000100110000001010100010110100101011001100010011001100101101001011100011000000110011001011100010110000101101001011010011001000110010001011010010110000101011001010010010001000011100,
	960'b000101000001011000011100000111100010000100100011001010010010100100101011001010110010101100101001001010010010100100101010001010100010110100101010001010010010101100101010001010000010100000101000001010010010101100101100001010110010101000101101001010010010101000101001001010010010100100101011001010110010101100101011001011010010100000101010001010100010110000101001001011010010101100101011001011000010101100101001001010000010100100101001001010100010110000101010001010110010101000101001001001110010100100100110001010000010100100101100001010110010101000101101001010000010100000101000001001100010011000101001001010110010100100101001001011000010101000101000001010010010100000101001001011000010110000101011001010110010100000101010001010010010100100101000001010100010101100101011001010100010101000100111001010000010100100101010001001110010101100101011001010110010101100101010001010000010101000101001001010100010100000101011001010110010101000100110001000000001111000011011,
	960'b000100000001010100011001000110110001111100100000000111110010011000101001001001100010010100101000001001100010001100100110001001010010001100101010001010010010010000100101001001100010001100100100001010000010010000100101001010100010100100100010001001010010011100100101001010000010011000100011001001110010101000101001001000110010011000100111001001000010100000100111001001000010101000101011001001100010010000100111001001110010010100100111001001000010001100101010001010100010010000100011001001100010010000100101001010000010010100100011001010100010101100100011001001010010011000100010001000110010011000100011001001000010101000101000001000100010011100100011001001010010100000100101001001000010100000101000001001000010011000100110001000110010010100100111001001010010011100101001001001110010010000101000001001110010010000101000001010000010001000101001001010010010010100100011001010000010010000100101001001110010011000100011001010000010011100011111000111100001111000010111,
};
localparam [0:85][959:0] b_picture = {
	960'b000110010001100100011010000111000010000000100001001000110010011100101001001010010010011000100101001001100010010100100111001001010010011100101011001010010010100000100011001000110010011000100101001001100010010100100111001010100010100000100110001000110010011100100100001000110010010100100100001001010010100100101001001001010010010000100101001000110010010000100100001001010010100000101000001001100010010000100001001001010010001100100100001001000010010100101000001001110010011100100110001001010010010100100011001001000010001000100101001010000010101100100111001001000010011100100011001000010010010000100001001001100010011100100111001001000010100000100110001001010010011000100101001001000010100100101010001001010010100000101000001001010010011000100110001001100010100000101100001010100010010000100101001001100010001100100101001001010010010100101001001010100010101000100010001000110010100000100100001001010010010100100101001010000010011100100011000111110001110000011010,
	960'b000110010001101100100000001000010010010000101101001011000010111000110101001100110011000100110100001100010010111100110001001100110010111000110011001101100011001000101111001100000010111000101101001100010011000100101100001100100011001000101111001011110011010000101110001011100011000100110000001011100011010100110101001011110011000100110001001011100010111100110010001100000011001000110101001100010010111100110000001011010010110000101111001100010010111100110010001100100010111100101111001100100010111100101011001011110010111100101101001100100011011000110001001100000010111100101001001010010011000000101111001100000011010000110010001011100011001100110000001100000011000100110011001100000011001000110100001011110011010000110011001100000011000000110010001100100010111000110100001101000010111000110010001100100010111000101110001100010011000000101100001100110011000100101111001100100010111100101110001011110011000100110001001011100010111100101001001001110010001000011111,
	960'b000111000010001000100101001011110010111000110001001110100011011000111011001110100011111100111001001110100011111100111010001110100011110100111010001111010011100100111110001110000011101101000000001110100011101100111011001101110011101000111000001110110011011000111010001110100011100000111110001110000011101100111010001110010011011000110110001110100011100100110111001110100011011100111101001101110011110100111000001101100011110000110111001110100011101100110011001101110011011000111100001110000011011000111000001101110011100000111011001101110011011100111000001110110011011100110111001101010011001000111001001101010011011100110101001110000011100100111100001111010011010100111010001111000011101000111010001110110011101100111000001111110011111100111001001111000011101000111011001110010011101100111001001110110100000000111101001110000011110100111011001110110011100000111100001110100011100100111101001110000011101000111101001101010011010100110010001011110010011100100011,
	960'b000111100010010100101100001110000011101000111010010000000100001100111111010000100100001101000011010001010100101001000101010000110100001101000011001111110100001101000011010000100100010101001011010001000100001101001010010001000100000101000100010000010100000101001000010010000100001001000010010001000011111001000010010010010100001101000011010001110100010101000010010000010100001000111110010000000100001101000010010000100100100001000010001111110100001101000000001110110011111001000010010000000100001001001001010000010011111001000100001111110011111001000011010000010100001101000101010001000100001001000000010000100011110000111100001111000100001101000111010010000100001101000000010000100100000000111111010000110100001001001000010010000100011101000111010000000100001000111111001111110100001001000000010001000100100101000110010001100100010001000111001111110100000101000010010000100100001101000111010001010100001001000011001111110011101100111101001101110011001000101100,
	960'b001000010010101100110101001110100100001101001000010000100100001101001011010001110100100001010000010100100101000001010100010100110100100101001000010010100100010101001000010101000101000101010000010101100100111101000111010010100100100001000010010010010101010001001111010011110101001101001001010001010100101001001100010010100100111001010010010011110101001101010100010010000100011101001000010001010100010101010000010011110100110101010010010011100100001101000100010010010100001101000101010100010100111101001010010100000100101101000101010001010100101101000111010010110101001001001111010100000101010101001011010001010100011101000110001111100100110101010001010011010101010001001010010001100100100001001000010001100100110001010011010100000101000101010111010011010100011001001001010010010100011001010001010101000100110001010001010101000100101001001000010011000100011101000111010100100101001101001011010100100100111101000110010001000100011000111111001110100011101100110011,
	960'b001001010010101000110110010000010100010001001001010010110100110101001101010100010101001001010001010100110101101001010100010100110101001101010000010011110100111101010001010101100101010001010101010101000100111101010001010100000100111101010001010011110101001101010110010101100101010001001101010100000100110101010000010100000100110101010001010110000101011001010100010011110100111101001110010100000100111101010011010100110101011101010101010100010100110101001110010011010101000101010001010100100101010101010110010100100100111001010001010011010100111101010011010100010101000001010101010101000101001101001101010011110100110101001110010011110100100101010111010110000101000001001111010101000100111101001101010101000101000001010000010110000101011101010010010100100101010001010000010100000101010001010010010100100101100001010101010100000101000101010010010100000101000101010101010011100100111101010111010100100100111101010001010011000100100001001000001111110011100100110100,
	960'b001010110010111000110111010010010100010101001001010101010101001001010100010101000101110001010011010101010110000001010110010110000101110101010110010110010101010001011010010100100101101001100010010100010101011001011011010100110101010001011001010110100101001001011100010111000101000001011010010101110101001101010010010111000101010101010011011000010101100101010010010110010101000101010100010101010101101001010010010101110110000001010100010100110101011101010010010100100101000001010110010011110101011101100000010100100101010001010111010100110101001001010111010101100100110001011101010111100100110101010110010101010101010101010100010100110101000101010111010111110101000001011001010101100101010101010010010110000101101101010010010110110101101001010110010111100101100001011011010101010101101101011000010100000101111101011001010100010101110001010100010110000101010001011101010110000101010001011011010101000101010101011001010011010101000101001010010010110011110000110111,
	960'b001010100011011000111011010000110100101001010110010101110101011101100010010110100101111001100000010110000101100101011010011001000101101001011101011001000101101101011101010111010101011001011010010110100110000001011001010111110110000001011000010111100101110101011010010110110101110101100001010110000110000001011100010111000110000101011000010110000101011001011101010111010101100001100011010110110101101101011111010101110101101001011011011000010101101101011100011000000101000101011010010110010100111101010110010110000101111001011000010111010101111101010110010110010101100001010111010101100101101101011100010100110110000001011110010101000101111001010110010110100110000101100001010101010110010001100100010101110101110101011110010110000101100101100001010111100101100101100101011000100101011101100000010111000101011101011100011000000101100101011011011001100101111101010111010111110101101101010111010110110110000001011001010110110101111101001111010011000100011100110111,
	960'b001001110011010101000001010000110101000001011000010110000110000001101001011001010101100001011101010111110101011001100001010111100101100101100011011000110110001001011100010111110101111101011010011000100101110001011001011010010110100101011011010110010110000101011101010111000110001101011110010111010110100001100101010110100101110101011111010101100101110001011111010110100110001001101000011000100101101101011011011000010101100101100001010111010101011001100101011001110101111001011000010110110101111001010101010111110101101001011000011001100110100101011101010101100110001001011001010101110110000101011000010110100110010101100001010101110110000001011011010110100101111101011110011000010110011101101000011000100101011101011111010101110101101001100000010111000101110101100001011000000110000001011001010111110101101001011100010110110101101101100010011010000110001001011100010110110110000101011001011000000101110101011011010111100101110001010001010010010100010000111101,
	960'b001100100011011100111101010010000100101101010111011001100110010001100110011001110110110001011101010110010101111001011101011001100110101001100010010111110110100101101001011000000101111001011111010110110110001101101100011001100110010001100111011001110101110101011110010111100101110101100101011010010110010001100010011010100101111101011001010111100101110001011110011010000110001101100001011001000110101101011110010110100101111001011001010111000110110001100100011000110110011001101010010111100101110001100000010110100101111001101001011000000110001101101001011001010101101101011011010110010101111101100101011000110110001001011100011000000101111101011101010111110101111001101000011010110110010001101000011011010110011101011101010111100110000001100011011011000110110001100011011001010110101101100111010111010110001001011010011000000110110001101001011000110110011001101100011001010101111101100101010111000110000101101011011000010101111001011000010101000100010000111010,
	960'b001100010011011100111101010010010100111001010101011000000110001101100110011001100110100001100000010111000110000001011101011000010110101101100110011001110110011101100101010111110101111001011100010111000110010001101011011000110110010001101010011001100101111001011101010111010101110001100111011011010110010001100011011010010101111101011010010111110101110101011101011010100110011001100101011000100110011001011101010111000101110101010111010111010110100101100100011000110110010101101010010111000101110101100001010111010101111101101001011000100110001101100110011000010101110001011011010111010101111001100000011000110110011001100000011000100110001001100000011000010110001101011101011001100110010101100111011001100101111001011101010111000110000101011101011000100110011101100110011001010110011001011101011000010101111001011100010111110110011001100111011001110110011001100111010111000101111001011110010111100101110101101000011000110101111001010111010100000100010000111101,
	960'b001010100011100001000011010010000101011001011011010110000110010101101110011010100110000001100011011000110101101101100011011001000101110001101011011010100110010101011111011001010110000101011111011001110110011001100110011101100111011001101100011001010110111101101000011010000110111101101100011011110111100101110110011010010110110101110001011010100110111001101100011001100111000101111000011101000110100001101101011011110110001101101101011010110110101001110101011101010111000001101000011011110110111101101001011011110110101001101001011101100111011001101101011010100110111101101011011010010110111001100111011010110111100101110100011001110111000101110000011011100111010101110001011010110111100001111000011010110110110001110000011010010110101001101110011010100110010001110001011011000101110101100110011010000101111001100101011010100110000101101000011011100110101101011010011001000110010001011101011000110110011001011100011010000110011001010110010011110100110000111111,
	960'b001011100011101101000001010010110100111101011101011000010101111001101000011000000101110101011100011000000110100101100000011010010110001001011110011010100101110101101001011011010110100101110111011111111001001010010111101000101010011110100011101001111010100010100100101000111010100110101000101000101010011110100100101001001010011110100010101000111010001110100110101001001010010010101011101000001010000010100100100111011001110110011100101000101001110110100001101000101001110010100000101000001001101010011010100111101010001010011100100111111010000010011100101000011001110010100000101001001010010010101000101000101010011010100010100111101010010010100101101001011010010010101010101001001010001110100101101001001010000010100010101010101010011010100001101000011001000110001011011110000111001001110100011000010110100101100100011000100110100101100000011010100101110101100101011001110101111001100010011000010110011001100100010110100101110101010100010101000100100001000000,
	960'b001011010011010100111111010101000101001001010101011000010110000001011100011000100110000101010110011001000111010101100001011000010110100001100011011001010110100001111010100000111001111010111010101111001011000110011100100011001000100010000101100000000111101101110110011100010110101001100101011000000110000001011111011000000101111101011101010111110110000001011101010111100101111101100010101011111011111010111100110000101100111011010010110110001101110111100000111000101110001011100011111000101110001011100010110111111101101111011000110100001100101111000010101110111011101110101010011000010101110001011101010111000101110101011111011000000101111101100000011000100110000001011111011000010110011001101110011101000111100001111011100001001000110110001010100100001010000110110101101110001011001010010110011111110111110101101110010111110110011001100100010110110110000001101001011000000110010001110000011000110101111101100100010110110101011101011001010011110100010001000011,
	960'b001010100011011101000100010011110101011001011100010101110101111001011010011000010101111101100101011011000110101001101100011010010110010101101100011110011001100010111000110001011010110001111011010100100011010100101110001011000010101100101010001010100010110000101110001011100010111000101110001011010010110100101011001011000010101100101001001010100010100100101001001010110010110000101010010100101010011010110010101110011100010111010001110110111110010111101010111100001111001111110011111100111111001111101111111010101110011011011101110100101100010110111010101101001010000001001001001010010010101100101101001100000010111100110000001011100010111100101111001011110010111000101101001011000010110100110001001011110010111100101110001011110011001000110011001100010011001100111111010110111000101010110101110000111010111010010101011111110110011101100001010111010101111101011111011001100110101001100111011010010110100101011101010101110101011101010100010010110100111001000011,
	960'b001010010011101001000111010010110101011101100001010101010101011001011111011000010101110101100110011010100110100101101101011011100111011010011010101111111011101010000111010011110011000000101110001100110011011100111010001110000011100000110111001101100011010100110111001101100011010100110100001101000011001000110010001101010011010100110100001101000011010100110100001101110011010100110011001011000100000101110011100100001001100110011110101000011010010010100110101010001010100110101010101010011010100110101000101001101010010110100010100111101001100110010001011100010011110000101111001101000011010100110110001101010011001100110011001101000011010100110101001101010011010100110110001100110011011100111001001111000100000001000001010000000011111100111110001111000011111000111111001101110011010000110111010110111001001111000011101101111000110001110011011001100101111101011100011001010110100101101000011011000110100001011101010110110101101101010101010011000100111001000010,
	960'b001011110011011001000000010100100100111101010001010111100110000001011101011001000110100001100001011001000111011001110011100011001011101110111010011100110011101100110001001101110011110000111111001111110011110100111100001111000011101000111101001111010011110100111101001111010011110100111100001110100011101000111001001111000011110100111011001111000011111000111110001111110011111000111100001111000011110100110111001101100011100000111000001110000011100000110111001101100011010100110100001101000011010100110101001101010011010100110110001101110011011100110111001110010011101000111011001110110011101100111100001111000011110000111100001111100011111100111110001111110100000001000000010000100100001000111101001111110011111001000000010000110100011001000101010001000100001101000011010000010100000100111101001110010011000001000011100000111011110110101001100000110110110101101001010111100110000101101110010111110101101001100110010111010101100101011000010100100100010101000001,
	960'b001011000011011000111110010011100100111101011000011001000101101101100010010111110110100101101000011010001000000110100011101111011000000100111000001011100011011000111010010000010100001101001000010101010110001101110010011111001000000010000010100000111000001110000001100000011000001110000011100000111000010010000100100001001000011110000111100010101000101110001100100011001000110110001101100011011000110110001101100011011000111010001110100011101000111010001110100011101000111010001110100011101000111010001101100011011000110110001101100011001000110010001100100011001000110110001101100011001000101110001001100001111000011110000110100001011000001110000011100000101000001010000011100001011000011010000110100010001000101010001011100010111000101010000110100000100111011101101000010110010100110101000100001111110011111000111000001011000100010010010011101110101001001001110110011010010110000101100011010111110110011101100101010111000101110101010011010101000100100000111101,
	960'b001010010011011101000010010010010101001101011110010111000110010001110001011001100101111001110001100001001010111010100111010011110010111100111011001111100011111101000110010110010111001110001100100111001010010010100101100111111001100110010101100100111001001110010001100100011000111010001100100011011000111110010000100100001000111010001111100100101001001010010010100100111001010010010101100101001001010010010101100101011001100010011000100110011001100110011001100110011001100010011000100110001001100010011000100110001001100110011001100110101001101010011011100110111001101110011010100110111001101010011011100110111001100010010111100110001001011110010110100101101001011010010111100101111001011110011010100110111001110010011100100111001001111010100010101010001010110010101001100111001000100001101110010101100100100001000011001111010011100100110001011000101011001010011101011101110110101001011011011001110110011101011011011001100110100001010111010011000100011101000000,
	960'b001011010011001101000000010010000101001001010101010111110110010101101011011010100110101001111101101101101000110001000001010000010100100101001011010011010101110101111111100111001010100110011110011111110101101101000000001100000010010100100011001001000010010000100100001001000010010000100100001000100010001000100011001000110010001100100011001000110010001100100011001001000010001100100011001001000010010000100100001001000010010000100011001000110010001100100011001000110010010000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100101001001010010010000100100001001000010010100100101001001010010010000100100001001000010010000100101001001000010010100100101001001010010010100101000001100000100001001100010100010001010001110100101100100110111001001011000010010110100100101000011001110000100101110100001101001000111100001100100011000010110000101101001011000110110000101011100010100000100001100111111,
	960'b001011110011011000111111010010110100111001011011011001110110010101101010011100001000111110110001011111000100010101010000010101010110001001100001011110111001110010101000100011000101010000101010000111000010001100101011001101010011101001000000010000010100000101000000010000000011111100111110001111000011101100111010001110010011100100111001001110010011100000111001001110000011100000111000001110000011100000111000001110010011100100111010001110100011101100111100001111010011111101000000010000000100000101000001010000000100000000111110001111000011110000111011001110100011101000111001001110010011100000111000001110000011100000111000001110000011100000111000001110000011100100111010001110100011101100111011001111000011111000111111010000000100000000111011001100110010101000011111000110110010110101011101100101001010001110001111011010100101100001011010010100110100100001000001100100011010011101111010011000100110011001110000011001000110001001011110010101010100011001000000,
	960'b001011000011010001000010010001110101001001010011010111010110100001110011100001101010111101110111010010110101111001101001011101110110111110001101101001111001011001001101000111110010001000110111010011010101101101100100011010110110101101101100011010010110101001101001011010010110100001100110011001100110010101100101011000110110001001100001011000000110000001100000010111110110000001100001011000000110000101100000011000100110001101100100011001010110011001101001011010010110100001101011011010010110100101101001011010100110100101101000011010010110100001100101011001000110001101100010011000100110000101100001011000010110000001100000011000000110000001100000011000010110000101100100011000110110010001100101011001110110100001101001011010010110101001101000011010010110010001011010010010010011010100100000001000010101100110011011100111000111101101011111011001100110010001010101010001011000111110100010011101110110001001100001011010010110011101011011010011100100100000111111,
	960'b001010000011100001000010010010000101001101011111010111000110100010000110101011010111111001001000011001010111111010001000011110011001010010100110011011010010010100100100010001000101101001100011011001100110011001100101011001000110001101100011011000100110001001100010011000100110000101100000010111110101111001011110010111010101110101011101010111000101101101011011010110110101101101011011010111010101111001011111010111110101110101011110010111110101111101100010011000100110000101100001011000100110000101100010011000100110001001100001011000100110000101011111010111010101111001011101010111110101111001011011010110110101101001011010010110110101101101011011010110110101110001011101010111010101110101011111011000000110000001100001011000010110001001100011011001010110011001101001011010100110011101011001001111110010000100101001011110111001111001111110011001010111000101110010010111100100011010010010100111100111011001011110011000000110000101010010010100110100110000111110,
	960'b001011010011011001000000010100100101010001010110011001000110110110100110100100010100110001100000100000101000111001111000100101011010000001001011000111100011110101011110011001110110001101100000011000000110000001011111011000100110010001100101011001000110010101100011011000110110001001100010011000110110001001100001011000000110000001100000011000000110000001100001011000000110000001100000010111110110000001100000010111110110000001100001011000100110001101100011011000110110001101100010011001000110010001100011011000110110001101100010011000110110001101100010011000010110000001100000010111110101111001011111010111110101111101011111011000000110000001100000011000000110000101100001011000010110001001100011011000110110001001100011011001000110010001100101011000100110000001100000011000000110001001100110011001100101101100111000000111110101101110011101100000000110010101111100011011010101001101000111100111101001000001101011010101110101010001010110010100100100001001000010,
	960'b001011100011011001000001010100010101000101010010011010011001010010100010010011000101100101111100100011110111011010010111100110100011110000101000010101000110100001100110011000000101110001011110011001000110011001100101011000110110001001100001011000000110000101011111011000000101111101011111010111100101110101011110011000000101111101011111010111100101111101011110010111100101111001011110010111100101111001011110010111100101111001011110010111110101111101011111010111110101111101011111011000000110000001100000010111110101111101011111011000000101111101011111011000000101111101011110010111110101111001011110010111100101110101011110010111100101111101011111010111110101111101011111011000000101111101011110010111110101111101100000011000000110000101100000011000100110010001100011011000110101111101011101011000010110100001100111010011100010001001001010100101100111101001100110011111100110001101001000010100111010010010000001010111110101010001011011010010100100011001000010,
	960'b001010010011110001000111010010100101100101100100011101101010110001011011010010100110010110001001011100101001001110011011001110010011000101100001011010110110010001100000011000000110001101100110011000010101101001011011010110110101101001011010010110110101101101011010010110100101101001011010010110010101100101011010010110010101100101011001010110000101100001011000010101110101100101011001010101110101011101011001010110100101101001011010010110100101101001011001010110010101101001011011010110100101101001011010010110100101101001011010010110110101101001011010010110100101101001011010010110100101101001011001010110010101101001011010010101110101100001010111010110000101100001011000010110100101101001011001010110100101101001011010010110100101101001011010010110010101100101011101011000110110011101100011010111100110000101101000011011100101110000101100010010011001001001101101011001000111001101010111001101110110111010100000011011000101110101010000010011000101000101000011,
	960'b001010110011100101000001010011100101001101100101100111011000001100111010010100000111010101101111100010111001111001000010001101100110011001101011011001000110000001100010011001100101110001011011010110110101101101011010010110100101100101011001010110100101101001011001010110010101101001011011010110110101101001011010010110010101100101011001010110010101100101011010010110010101100101011010010110100101100101011001010110100101100101011010010110100101101001011011010110100101101001011011010110110101101001011011010110100101110001011011010110100101101001011010010110010101100101011001010110010101100101011001010110010101101001011010010110100101100101011001010110010101101001011010010110100101101101011011010110110101101101011011010110010101100101011001010110010101101001011010010110100101110001100010011001110101111101100001011001110110111001100100001010110101001110000110010111110110001001100000010001000011010010010111100010000101101101011000010011000100011101000001,
	960'b001011110011010100111111010101010101010101111000101010100100000000111111010111110110011001111100100111100101101000110011011010110110110001100110011000000110010101100011010110110101101001011011010110100101101101011100010110110101101101011011010110100101100101011011010110110101101001011011010110100101101001011010010110100101101001011010010110010101101001011001010110010101101001011010010110100101101001011010010110010101101001011010010110010101101001011001010110100101101001011010010110100101101001011011010111000101101101011010010110100101101001011010010110100101101001011001010110100101101001011011010110100101101001011001010110100101101001011010010110010101100101011001010110100101100101011010010110100101101001011011010110110101101101011011010110110101101001011010010110100101101101011010010111010110100101100101011000110110011101101101011001010010111001100101011110000101010101011100010010010011000001010000101000010110101101010001010100010100001000111111,
	960'b001010100011100001000001010010000101101110100001011101010011000001000010010101110110110110010110011111010010111101100101011011100110010001100001011010100110001001011110010111010101110001011100010110010101100101011010010110110101101001011010010110010101101001011011010110100101101001011010010110100101101001011001010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110010101100101011010010110100101100101011010010110100101101101011011010110010101100101011010010110100101101001011010010110100101100101011001010110100101101001011010010110100101101001011011010110010101100101011010010110100101100101011010010110010101100101011010010110010101101001011010010110110101101101011011010110110101101001011011010110010101101001011011010111000101111101101001011001100110010001101000011011110101111100101110011110010110010101001110010010010011011000100111100011011001000001010110010011110100110100111011,
	960'b001010100011011001000010010001100111001010101011001110110011000100111110010100011000010110010011001110010101100001110000011010000110001101101000011000110101110001011110010111000101101001011010010110000101100001011001010110110101101001011010010110100101100101011010010110100101100101011010010110100101101001011010010110100101101001011010010110100101100101011010010110100101101001011001010110100101101001011010010110100101101001011010010110110101101001011001010110100101101001011010010110100101101001011001010110100101101001011001010110100101101001011001010110010101101001011010010110100101100101011001010110100101100101011010010110100101101001011001010110100101101001011010010110010101100101011001010110100101101001011010010110100101101001011010010110100101101001011010010110010101101001011011010110110101110101100000011010000110010101100110011010010111000001001101010001100111011101010001010001010011011000100110010011101010100101101010010010100100001100111110,
	960'b001100100011100000111011010100101000111110000001001001110011000000111110011010011001001001100011010000010111000001101001011001010110100101100110010111010101110101011111010111010101101101011010010110100101101001011010010110010101100101011010010110110101101001011001010110100101101001011010010110100101101001011010010110100101101001011010010110010101100101011010010110010101101001011010010110100101100101011010010110010101101001011001010110100101101001011010010110010101100101011010010110100101100101011001010110100101101001011001010110100101101001011010010110010101101001011010010110010101100101011010010110100101100101011001010110100101100101011001010110100101100101011010010110010101100101011010010110010101101001011010010110100101101001011010010110100101101101011010010110100101101101011100010111010101110101011111010111110110101101100011011001010110101101101111001110000110010001100010010001110011100100101100001001011001100010000011010101010100010000111110,
	960'b001100000011010100111100010111111010010001001010001010000010111001000101011111011000101000111101011010000110110101100110011000100110101101011111010111010101110101011101010111000101101101011010010110110101101001011010010110100101101001011010010110010101100001011010010110100101101001011010010110100101101001011001010110010101101001011010010110100101101001011010010110010101101001011011010110010101101001011001010110100101101001011001010110100101101001011001010110010101101001011010010110010101101001011010010110100101101001011010010110100101101001011010010110010101101001011001010110100101101001011010010110010101101001011010010110100101101001011010010110100101100101011010010110110101101001011010010110100101100101011010010110010101101001011010010110100101100101011011010110100101101001011100010111000101110001011101010111010110001001101000011000110110100001101110010111100100000101101110010011010011101000101101000111010110100010011011010110010100010000111111,
	960'b001010000011010101000011011100011001101100101100001010010011000001010111100001000110010101001001011100000110100001100010011001110110000001011110010111010101110101011011010110010101100101011001010110100101101001011010010110100101101001011010010110100101101001011001010110010101101001011010010110010101101001011001010110100101101001011001010110010101101001011010010110100101100101011001010110010101101001011010010110100101100101011001010110010101100001011001010110010101100101011001010110000101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011010010110010101100101011010010110010101100101011010010110010101100101011010010110010101101001011010010110100101101001011010010110010101101001011010010110110101101001011010010110010101101001011011010111000101110001011101010111010101110101100101011001010110001101101001011100010100001101100010010101110011111000101111001001100011100110011110011000110100101100111110,
	960'b001010100011011001000101100010100111100100100001001010010011100001100111100000010100100001100110011010000110010001100001011001010101101001011110010111100101110001011010010110010101100001011001010110100101101101011010010110100101101001011010010110100101101001011010010110100101101001011010010110110101101001011001010110100101101001011001010110100101101001011001010110100101100101011000010110010101100101011001010110000101100101011001010110000101100001011001010110000101100101011000010110010101100001011001010110010101100101011001010110000101100101011000010110010101100001011000010110010101100101011001010110100101100101011010010110100101101001011001010110010101101001011010010110100101100101011010010110100101100101011010010110100101100101011010010110100101101001011010010110100101101001011011010111000101110101011101010111000101110101011100011010000110000101100101011010100101111001001101010111010100010100110001001010010010000010010000011111000100100100111111,
	960'b001011010011000101001100101000010101001000100100001010010100001001101100011100010100101101101101011001000101111001100110011000000101110001011101010111010101110001011011010110110101100101011010010110010101101001011010010110100101100101011001010110100101101001011010010110010101100101011010010110100101100101011001010110010101100101011010010110100101101001011000010110000101100101011001010110010101100001011000010110010101100001011001010110010101100101011000010110000101100101011001010110010101100001011001010110010101100001011001010110010101100001011000010110010101100101011000010110010101100101011001010110010101100101011000010110010101101001011010010110100101100101011010010110100101100101011001010110100101101001011001010110010101101001011010010110100101101001011010010110100101101001011011010110100101101001011101010111000101110001011001011000110110000101100000011001000110101101001000010111110100100100110111001010110001100101101110100010100100101001000010,
	960'b001010100011010001011101100111100011011000100110001011010100110001101101010111100101100101100111011000010101111101100101010110100101101101011100010111000101110001011100010110110101101001011010010110110101101001011010010110100101101001011010010110100101100101011010010110100101101001011010010110100101101001011010010110110101100101011001010110010101100101011001010110000101100001011001010110000101100101011001010110000101100101011001010110010101100001011001010110010101100001011000010110010101100101011001010110000101100101011001010110010101100001011000010110000101100101011001010110010101100001011000010110010101100001011001010110000101100101011010010110100101101001011001010110010101101001011010010110010101101001011010010110010101100101011010010110100101101001011010010110100101101001011011010101110101011101011100010111010101110101011100010111100110010001011110011000100110110001010010010110100100111000111100001010100001110101001010100101000101101000111111,
	960'b001001110011101001101111100011110010010100100111001100110101000001101001010101100110001101100101010111100110001001100000010110100101101101011101010111000101100101011010010110110101101101011010010110110101101101011010010110100101100101011001010110010101100101011010010110100101100101011010010110100101100101011010010110100101100101011001010110010101100101011001010110010101100101011000010110000101100101011000010110010101100101011001010110010101100101011001010110000101100101011000010110010101100001011000010110010101100101011001010110000101100101011001010110010101100001011001010110000101100101011000010110010101100001011001010110010101100101011000010110100101101001011010010110100101100101011001010110010101101001011001010110100101100101011001010110100101101001011010010110110101101101011011010110010101101001011011010110110101110001011101010110100110010101011101010111110110011101100000010101000101001100111111001011010010001000101111100101100110001001000010,
	960'b001010100011100001110111011110110001111100101000001110010101001001100111010101010110011101100100010111000110010101011110010111000101101101011011010110110101101001011011010110100101101001011010010110100101101001011011010110100101101001011010010110100101101001011001010110100101101001011001010110100101100101011001010110100101100101011000010110000101100101011001010110100101100101011000010110010101100101011001010110010101100101011001010110010101100101011000010110100101101001011001010110010101100101011000010110000101011101011000010110000101101001011010010110010101100001011001010110000101100101011001010110010101100001011001010101110101100101011000010110100101101001011010010110100101101101011001010110010101101001011001010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011011010110110101110001011100010110010110001001011110010111100110001101100111010101010101011001000100001100100010011100100001100010110110010001000010,
	960'b001011010011110101111110011000100010000000101011001111100101001101100100010111010110100101100010010111000110010101011011010110110101101101011010010110010101101001011001010110100101100101011001010110100101101001011010010110100101101001011001010110100101101001011010010110010101101001011010010110100101101001011001010110100101100001011000010110010101100101011001010110000101100001011001010110000101100001011001010110010101100001011001010110010101100001011001010110010101101001011001010110010101100101011001010110000101100101011010010110010101100001011000010110010101100001011001010110000101100001011000010110010101100101011001010110010101100101011010010110100101101001011010010110100101101001011001010110010101101001011010010110010101101001011010010110100101101001011010010110100101101001011011010110100101101101011010010110110101101101011100010110100101111001100011010111010110000101101000010111000101011101000101001101000010100100011100011111000110110101000000,
	960'b001010010100001010000100010011110010001100101111001111100101000001011111011000100110100001100001010111010110001001011010010110110101101101011011010110110101101001011000010110110101101101011010010110110101101001011011010110100101101101011010010110100101101001011010010110010101100101011010010110100101101101011001010110010101100101011001010110000101100101011001010110000101100001011001010110010101100001011001010110100101100001011000010110000101100001011000010110000101100101011000010110010101101001011000010110010101100001011010010110010101100101011001010110000101100001011000010110000101100101011001010110010101100101011001010110000101100101011001010110100101101001011001010110010101100101011001010110010101100101011010010110010101101001011001010110010101101001011010010110100101100101011010010110110101101001011010010110110101101101011011010111000101111101100101010111010110000101101001011000010101101001000100001110000010100100011010011011110111010101000000,
	960'b001010110100000110000110010001010010010100110011010000010100110001011110011001110110100001100001010111110110001001011010010111000101110001011100010110110101101001011000010110100101101001011010010110100101101001011010010110100101101001011010010110100101100101011010010110010101101001011010010110010101101001011011010110010101101001011000010101110101100001011010010110000101100001011001010110000101100101011000010110010101100001011001010110010101100001011000010110010101100101011000010110000101100101011000010110010101101001011000010110010101101101011001010110010101100101011001010110010101100101011010010110100101100001011001010110100101100001011000010110100101101001011001010110100101101001011001010110100101101001011010010110010101100101011001010110100101100101011010010110100101101001011010010110100101101001011010010111000101101101011101010111000101111101100100010111110110001001101001011001010101110101000110001110110010110000011001011001110111011000111110,
	960'b001011110100011110000110010000000010010100110100010001000100100101011111011010110110100101100011010111110110010001011011010111000101110101011100010111000101101101011010010110100101101101011010010110010101101001011010010110010101100101011010010110100101101001011010010110010101100101011010010110010101101001011001010110010101100001011001010110000101100101011000010110010101100101011000010110010101100001011001010110010101100001011001010110000101100101011000010110000101100101011000010110000101100001011001010110010101100001011000010110010101100101011000010110000101100101011001010110010101100001011000010110000101100101010111010110000101100101011010010110010101101001011001010110100101100101011001010110010101100101011010010110010101101001011010010110010101101001011010010110100101101101011001010110100101101101011011010110110101101101011010010111000101110101100101010111110110010101101000011011100101110001000110001111100010111100011010011001010111101001000000,
	960'b001010110100000110000111010000100010100000111001010001010100011001100001011100010110101101100101011000010110011101011100010111000101101101011100010110110101110001011010010110100101101001011010010110100101101101011010010110100101100101011010010110100101101001011001010110010101101001011001010110000101101001011010010110100101101001011001010110000101100101011001010110000101100001011001010110010101100101011001010110010101100001011001010110010101100101011001010110010101100001011000010110010101100101011001010110010101100001011001010110010101100001011000010110010101100001011000010110010101100101011000010110000101100101011000010110000101100101011010010110100101101001011001010110010101101001011001010110100101101001011010010110010101101001011010010110010101101101011010010110100101101001011010010110100101101001011100010111000101110101011100010111000101110101100111011000100110011101101100011100110101111001000101010000100011001000011110011001010111101101000010,
	960'b001001010100001110001000010001010010101000111011010010000100010001011110011101010110110101100111011000100110100001011101010111100101110001011100010110110101101101011011010110100101101001011011010110110101101001011010010110100101100101011001010110100101100101011010010110100101100101011001010110100101101001011010010110110101100101011010010110010101100001011001010110000101100001011001010110010101100101011001010110000101100001011001010110010101100001011010010110010101100001011001010110010101100101011001010110000101100101011001010110100101100001011000010110000101100001011001010110000101100001011000010101110101101001011010010110010101100101011010010110010101100101011010010110100101101001011010010110100101101001011001010110010101101001011010010110100101101101011001010110100101101101011011010110000101101101011100010111000101111001011101010111110110000001100110011000100110100101101111011101000101101001000101010001010011010100100001011010010111111000111111,
	960'b001010010011111010000100010001110010101100111101010100000100001101010111011101010110111101101000011001000110100101011111010111110101110001011011010111000101110001011100010110110101101101011001010110100101101001011010010110100101101001011010010110010101100101011010010110010101100101011010010110100101101001011010010110010101100101011010010110110101100101011010010110100101101001011000010110000101100101011000010110000101100101011001010110000101100101011010010110010101100101011001010110100101100101011001010110100101100101011001010110010101101001011001010110000101100001011000010110000101100101011001010110100101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110010101101001011010010110100101100101011010010110110101101001011010010110110101101101011010010110000101110001011011010111000101111001011110011000000110001101101000011000110110101001110001011101010101011101000101010010100011100000100000011010000111011101000100,
	960'b001010010011111110000100010010010010110001000001010101000100001001010001011101100111010001101010011001000110100101100001010111110101110001011110010111010101110001011100010110010101101001011011010110100101101001011011010110100101101001011010010110010101100101011011010110010101100101011010010110110101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110010101100101011010010110100101100101011010010110010101101001011001010110010101100101011001010110010101100101011010010110010101101001011001010110010101101001011001010110010101101001011010010110010101100101011010010110100101100101011001010110010101100101011010010110010101100101011010010110100101100101011001010110100101100101011010010110010101101001011011010110100101100101011010010110100101101001011010010110110101110001011011010111010101111001011110010111110110011001100111011001100110110001110101011101110101000101000100010100110011100100100000011010100111100001000011,
	960'b001001110100000010000110010011000010111101000110010111110100010001001010011101000111011001101101011001110110100101100110010111110101110101011111010111100101110001011101010110010101101101011011010110100101101001011011010110100101101001011010010110100101101001011001010110100101101001011001010110100101101001011010010110010101100101011010010110100101101001011001010110010101101001011010010110100101101001011010010110100101101101011010010110010101101001011010010110110101101001011011010110100101101101011010010110100101101001011011010110100101101001011010010110100101101001011010010110100101101001011010010110010101101001011010010110100101100101011010010110100101101001011010010110010101101001011010010110100101100101011010010110010101101001011010010110010101101001011010010110110101101001011011010111000101110001011011010111000101111001011111011000010110101001100101011010010110111001110110011101000100101001001100010111000011110100100101011011110111101101000010,
	960'b001010000011110010000000010100110011001101001100011010000100100101000100011010100111110001101111011010110110100001101010011000010101111101011110010111010101110001011100010110100101101001011011010110100101101001011010010110100101101001011010010110100101101001011001010110100101101001011010010110100101101001011001010110010101101001011001010110100101101001011010010110010101101001011010010110100101101101011010010110110101101001011010010110110101101101011010010110110101110001011100010110110101101101011010010110110101101101011011010110110101101001011011010110110101101001011010010110100101101001011010010110100101101001011011010110100101101001011010010110100101101001011010010110100101101001011001010110100101101001011010010110010101101001011011010110100101101001011010010110100101101001011001010111000101110001011101010111100101111001100000011000110110110101100110011010010111000101111101011010010100010001011011011010000100001100101010011101000111001101000011,
	960'b001010110011101001111001010111100011101101010101011100100101111000111101010110100111110101110100011010110110100001101101011000100110000101011110010111000101110001011100010110110101101001011011010110100101100101011010010110100101101001011010010110110101100101011010010110100101101001011001010110100101101001011010010110100101100101011010010110100101101101011011010110110101101101011010010110100101101101011011010110110101101001011011010110110101101101011100010111000101101001011010010111000101101101011011010111000101101101011011010110110101110001011011010110110101101101011011010110100101101101011011010110110101101001011010010110100101101001011010010110010101101001011001010110010101101101011010010110010101100101011010010110010101101001011010010110100101101001011010010110100101101101011001010111000101110101011111010111110101111101100000011001100110101101101000011010110111011101111111010110000100000001110010011011100100010100110000011111000110011001000011,
	960'b001010100011101001110001011001010100000001011100011101000111101100111011010011000111101101111001011011000110011101101100011001100110000001011111010110110101101101011100010111000101101001011011010110100101101001011010010110100101101001011010010110100101101001011010010110100101100101011010010110010101101001011010010110100101100101011010010110110101101001011010010110110101101101011010010110110101101101011011010110110101110001011100010111000101110001011101010110110101101101011011010111010101110101011101010111000101110101011101010111000101110001011100010111000101110001011011010110110101101101011011010110100101101001011011010110110101101001011010010110110101101001011010010110010101100101011010010110010101100101011010010110100101101001011010010110100101101001011010010110100101101101011010010111000101110101011101010111010101111101100001011010100110011101101001011100000111110001110110010010000100011010001011011011110100011100110101100001100110001000110100,
	960'b001010100011100001101001011101100011111101011111011100111000111001001010010000100110101001111110011100010110100101100111011010100110000001011110010110110101110001011100010111000101101101011011010110110101101001011010010110100101101001011010010110100101100101011010010110100101101001011010010110100101100101011010010110100101101001011010010110100101101001011010010110100101101101011010010110110101101101011100010111000101110101011101010110110101110001011101010111010101111001011110010111010101111001011110010111010101111001011101010111100101111001011101010111010101110101011100010111000101110001011100010111000101101101011010010110110101101001011011010110100101101001011010010110100101100101011010010110100101101001011011010110100101101001011010010110100101101001011010010110100101101101011011010110110101101101011100010111010101111101100100011010110110011101101011011101000111111101100001001111110101111110010000011010110100111000111011100010110101100100111011,
	960'b001100010011010101010111100001100011011001100011011100101001001101101010001110000101001101111101011101110110110001100110011010100110011001011100010111000101110001011100010111000101101001011011010110110101101101011010010110100101101001011011010110100101101001011011010110100101101001011010010110100101101001011001010110100101101101011011010110110101101101011010010110110101110001011100010111010101110001011100010111000101110001011100010111000101110001011110010111110101111101011111010111110101111001011110010111100101111101011111010111010101110101011111010111100101110101011100010111000101110001011100010110110101110001011100010110110101101001011010010110100101101101011010010110110101101101011010010110100101101001011010010110100101101001011010010110100101100101011001010110110101101001011011010111000101101101011100010111100101111001101011011001110110100101101110011110010111101001001101001111001000100010001101011010000100111101000011100011010100110100111010,
	960'b001100010011011101001011100010110011011001011100011011011000011110001111001111010100010001101110011110100111000001101001011001000110101001100000010111010101110001011010010111000101101101011011010110100101101001011011010110100101101101011011010110100101101101011011010110110101101101011011010110100101101001011011010110110101101001011010010110100101101001011011010111000101110001011100010111010101110101011011010111000101110101011101010111000101110101011101010111010101110101011110010111100101111001011110010111110101110101011110010111100101111001011110010111100101110101011100010111010101110001011100010110110101110101011101010111000101110001011011010110110101101101011011010110110101101101011011010110110101101001011011010111000101101101011011010110110101101001011001010110110101101101011100010110110101101001011101010111010110011001101000011001010110101001110000011110110110000100111110010100011001011101111100010111110011110101011101100000000100100100111101,
	960'b001010100011010101000111100000100101000000111110011001110111100010010111011000110011101001010011011110000111010101101100011001100110001101101001010111010101101001011010010111010101110001011011010111000101110001011100010110110101101101011011010110110101101101011011010110110101101001011011010110100101101101011011010110100101100101011010010111000101110001011101010111010101110101011101010111000101110001011101010111010101110101011101010111000101110101011100010111010101110101011101010111010101111001100000010111110101111001011101010111110101111001011101010111000101110101011101010111010101110101011101010111000101111001011101010111010101110001011100010110110101100101011001010110110101101101011011010110110101101001011011010110100101101101011100010111000101110101011100010111000101110001011100010111000101110101011101011000010110100001100001011001010110101101110110011100110100011100111010011110001000000001101000010111000010010001111101011100010100101100111111,
	960'b001010110011101101000100011100010111100100011011010111110110011010000100100011000011111001000001011000110111100001110000011010000110000101100001011001110101101001011010010111000101110001011100010111000101101101011100010111010101101101011100010110110101101101011011010110110101101001011010010110100101101001011011010110110101101001011011010111000101110001011011010111010101110101011110010111010101111101011100010111010101110101011110010111100101111101011111011000000110000001011111010111110110000001100001010111110110000001100000010111110101111101100000010111110101111101011110010111100101111001011110010111000101111001011101010111000101110001011100010110110101101001011010010110100101101001011010010110100101101001011011010110110101101101011011010111000101110001011101010111000101110001011010010111000101110001100000011001110110000001100011011010010111000101111001010110000011111001001100011111100110011001010100010010010010010010010100011001010100100000111111,
	960'b001011110011010101000001011001011001001000100101001111010101001101100001011111110110000100111001010001110110110101110011011010110110010001100001011000010110010101011100010110110101101001011010010111010101110101011110010111100101110101011101010111000101110001011100010111000101110001011100010111000101101101011100010111010101110001011100010111000101111001011011010110100101110001011101010111000101111001011110011000000101111101100000011000010110000101100001011000100110000101100010011000100110001001100010011000100110001001100010011000010110000101100000011000000110000101100000010111100101111001011110010111100101111001011110010111010101110101011101010111010101110001011100010110110101110001011011010111000101110001011100010111000101110001011100010111010101111001100000010111100101110101011100010110110110000001100111010111110110001001100101011011000111100001100100010000110011101001100101011000010100111001001111001000010101010110001110010101010100001101000100,
	960'b001010110011010101000010010110001000011101100000000100000100110101001011010110110111001101000110001111010101000001110000011011110110011101100011010111010110000001100111010111110101100101011100010111000101110101011110010111100101111101011110010111010101110101011101010111010101111001011110010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011110010111100101111101100000011000000110001001100011011000100110001101100100011000110110001001100100011001000110001101100100011000110110001101100100011000110110001101100011011000110110010001100001011000100110000101011111011000000101111101011110010111010101110101011110010111100101111001011101010111010101110101011101010111010101110001011100010111010101110101011101010111010101111001011111010111000101110001011101011000110110010101011110011000010110010001101010011100110110101001000111001110110100110001010101010001100100000000111110000011101000100101110101010011110100111001000100,
	960'b001010000011100101000110010011010111001110010101000101010010101101000110010010000101001101011100001110110100000001011000011100000110101101100110011000100101110101011101011001010110010001100000010110110101101101011100010111100101111001011110010111110101111101011111010111100101111001011100010111000101110001011011010110110101101101011100010111000101110001011101010111110101111101100000011000010110000101100010011000100110001101100001011001000110010001100100011001000110001101100100011001000110010001100101011001010110010001100100011001000110010001100101011001000110001101100010011000100110001001100001011000010110000001100000010111110101111001011101010111010101110101011100010111100101110101100000011000010101111001011110010111110101111101011111010111100101111001011101010111010110010001101000011001000101111001100001011000110110011101110001011011100100101100111110001111110100111000111100001101110100000000010100001111101001100101011110010011000100111101000011,
	960'b001010110011011001000010010100110101100110001111010100110000010000111100001110100100001001001100010100100011101001000000010111010110111101101100011001100110010001100000010111010110000001100110011001110110001001100001011000000110000001100000011000010110000001100001011000000101111101011110010111010101110001011101010111010101110001011100010111100101111001011111011000000101111101100001011000010110001001100010011000100110001101100011011001000110010001100100011001010110010001100100011001010110010101100101011001010110011001100101011001000110010101100100011001000110001101100011011001000110010001100010011000010110000001100001011000000101111001011111010111100101111101011110010111100101111101100000011000000110000001100000011000000110000001100011011001000110010101100110011010000110100101100011011000100110010001100101011010100111000001101101010011010011111000111011010001010011010100110001001100100010100100001000100000100111111101011100010011110100010001000010,
	960'b001011000011011000111111010011110101000101110101100101010001101000010101001111000011100000111111010010000100100100111000010000000101101001110010011011000110101101100111011001010110010101100001011001000110101001101011011010110110101101101010011010100110101101101100011010110110101101101000011010000110100001101010011010100110100001100111011010000110100101101010011010110110101001101010011010100110101001101010011010110110101001101011011011000110110001101100011011000110110001101110011011010110110001101101011011010110110001101100011011010110110101101100011011000110110001101011011011000110101101101011011010110110100101101000011010100110100101101001011010000110100001101000011001110110100101101000011010100110110001101101011010100110101101101010011010110110100101100111011001010110010101100110011001110110100101101101011100010110101001001001001111100011100000111101001100100010111000101010001011100000010001000101100110010110011101010101010101100100011100111110,
	960'b001010000011100101000001010010000101001001100110100100010110011100000001001000010011011000111001001111110100000101000100001101110011110001010100011101010111010001101011011011000110101001101001011010010110100001100111011001110110100101101000011010010110100001100111011001110110011101100110011001110110011001100110011001100110010101100101011001100110011101100110011001110110011001100111011001100110100001100111011001110110011101101001011010000110100101101001011010010110101001101010011010100110101001101001011010010110100101101010011010010110100001101001011010010110100001100111011010010110100001100111011001100110011101100111011010000110011101100101011001010110011001100110011001100110011001100110011001110110011101101001011001110110100001101000011001110110011101101000011010110110110001101010011011110111001001110100011000110100100000111110001101000011010100110000001011110010011000101101000011010001001110001011100001100110100101010010010011100100101000111111,
	960'b001011000011001101000001010001110101001101011001011101001001111100110011000000000010100000110101001101110011101000111101010000110011101000111000010001110110101101111011011101110111000101110000011100010110111001101101011011000110110101101110011011010110110101101100011011000110110101101011011011000110101101101011011010100110101001101010011010110110110001101011011011000110101101101011011010110110101101101011011011010110111001101110011011110110111001101101011011100110111101101111011011010110111001101111011011110110111001101110011011110110111101101111011011110110111001101111011011010110110001101011011010110110101101101011011010110110101101101011011010110110101101101011011010100110101101101010011010110110110001101100011011010110111101101111011100100111000101110001011100100111001101111000011101110110111101010100010000110011110000110110001100110010110000101100001001000010100100010100000000110110011010011011011011010110001101011110010010110100010000111111,
	960'b001011110011010100111110010011000100110101011010011011001000101010001111000100110000010100101010001101010011010100111010001111000100100101000101001110010011110101010010011101011000100010000010011110110111100001110111011101110111011101111000011110000111100001110111011101100111011001110011011100110111000101110000011100000111000001101111011100000111000101110010011101000111000101110010011100100111001101110100011101010111010001110101011101010111010101110100011101010111011101110111011101010111010101110111011101110111011001110101011110000111011101110110011101100111011101110111011101010111010101110011011101000111001101110010011100100111000101110001011100010111001001110010011100010111001101110010011101000111010101110111011101110111100001111000011110110111110101111110011111010111110001110011010111100100100100111101001110000011101000110011001011000010100100100011001010100001011000000010001111011010000101111101011001000110000001100000010101010100011001000000,
	960'b001010110011010101000001010010100101000101010011011000110111000010011010011101000000011100000110001011000011100000110010001101110011101001000111010101100100100000111011001111100100111001101100011111111000100010001001100010011000100110001010100010111000101010001001100010001000011010000101100001001000001010000010100000011000000010000000100000011000000110000000100000011000001010000100100001011000010110000111100001101000010110000101100001011000011010000110100001101000010010000100100001001000010110000101100001001000010110000101100001111000011110000100100001001000011110000110100001101000011010000110100001011000001110000100100001001000001010000011100000101000000110000010100000011000001110000100100001101000010110000111100001111000100010000110100001101000010101111011011011000101100001000111001111100011101101000001010000000011000100101011001001100010010000101111000101110000001100100001100101111000000101101010011010000110010001011010010011010100100001000001,
	960'b001010000011100101000011010001110101011001011111010101100110100101111010100111010101110100000011000001100010010100111011001011100011001100110110001111010101000001011010010011000011111100111010001111100100101101010111011001010110110001110010011101010111011001111000011110100111110001111110100000011000001010000100100001011000011110001001100010111000110010001011100011001000111010010000100100001001000010010010100100111001010010010101100101001001010110010110100101101001011110011000100110011001100110011000100110001001100010011000100110001001100010011000100110001001011110010110100101011001010010010010100100011000111110001110100011001000101010000111100001011000000101111111011110110111100101111001011110000111001101110001011100000110110101100101010110110101000101000101001111110011110000111110010001010100100000111100001011110010101000100110001010010011000000010101000001000001011010000110100100000110111101011100011001000110001001010001010100110100101100111110,
	960'b001011100011100101000001010011110101001101011011011000000101110001100100011101011010001101010011000001100000010100011001001110100011000100101101001100100011011000111110010010110101001101010101010011110100011001000011010000010100000101000011010000110100010001000111010010010100100001001001010011000100110101001101010011100100111101010001010100110101010101011000010110010101101001011011010110100101101101011100010110110101110101011101010111110110000001100010011000100110001001100011011000110110001101100010011000100110000101100010011000110110001101100010011000010110000101011111010111010101101101011010010110010101100001010110010100110101000101010010010100000100110001001010010010100100100101001000010001100100010001000011010000100100000101000010010000010100001001000110010001010100011001000110001111000011001100101101001001110010010000110001001011100000111100000101000100100111111110011101011010010110011001100011010101110101010101010110010100100100010001000000,
	960'b001011010011011101000010010101000101000001010001011000110110001001011110011010100111110010011110010101100000011000000101000010110010110100111001001011010010110000110100001100100011011000111011010001110101001001010000010011100100111001001101010011010100110001001100010010110100011101000011010000110100001001000010010000100100000001000000010001000100011101001010010011000100110101010000010100110101010001010011010101010101100101011011010111110110000101100010011000100110001101100011011000110110010001100001011000010101111001011111010111110101110001011011010110010101011101010010010011010100101101001011010010000100011001000101010010000100100001001000010010000100100001001000010011000100110101001101010011110100111101001110010011100100111001001111010100100100101101000010001111000011010000110000001011100010110000101001001011100011010000011110000010000000010100010111011111101001100001110111011000110101111001100011010110100101011001011010010010110100010001000010,
	960'b001010100011101101000110010011000101011101011010010110010101110101011110010111110110001110000000101001010110011100001111000001000000011100010100001100000011101000110001001010010010101100110000001100010011010100110010001100110011010000110011001101000011010000110011001100010010111100101101001011010010110100101111001011100010110000101010001011000010110100101101001100000011000100110000001100100011001000110011001101010011100000111001001110010011101000111010001111000011110000111100001111010011111000111110001111100011110100111100001110100011100000111010001110000011010100110011001100010011000000110001001011110010110100101011001010110010101100101101001011010010110100101110001011000010111000110001001100110011011000110111001110000011011100110100001101000011000100101110001011110010110000101011001011010011011100111001001001110000110000000110000001000010001010001001100111110111011101100111011011100110001101011011010111010101100101010000010011100101000001000111,
	960'b001010110011101001000100010011000101010001011001010110010101110001011010011000100101111101101010011110001010000110000001001000110000011000001001000010000001101000111001010001110011111000110000001001110010011100101001001010110010101100101101001011100010111100101110001011000010110100101100001011000010101100101100001010110010100100101001001010000010100000101001001011000010110000101100001011000010110100101111001100000011000100110000001100000011001000110100001101000011001100110011001101010011010100110011001101000011010000110011001100100011000100110010001100010010111000101101001011010010110000101010001010100010101100101011001011010010110100101011001010100010100100101001001010100010110000101011001010100010101100101011001011010010110100101100001011000010101100101011001100000011101101000100001111110010101100001111000001000000010100000110001111111001011110001101011011110110011101100110011001000101111001100000010110110101010101010110010011010100100101000010,
	960'b001011110011010101000000010101010101000001010010011000000101111001011100011000100110011001011100011010000111110110010000100110000100111000001110000001010000011100001011000111110100011101100011011001100101101101010010010100000101000001010001010011110101000001001111010011100100111001001111010011010100110001001010010010010100011101000110010010000100100001000111010010000100100001000111010010010100100101001011010010110100101001001001010011010100111001010000010100010101000101010001010100010101001001010010010100010101000101010001010011100100110101001011010010100100100101001000010010000100011001000101010001000100010101000100010000110100010001000101010001010100100001000111010001110100011001000110010010000100100001000111010010010100100101001000010010100101000101011010010110100100010100100110000011110000010100000111000001100001110001101010101000001000001001101110010110100101111101101010010110100101111101100101010110010101010001010011010100000100000101000010,
	960'b001011100011100001000000010010100100101101011000010111100101111101100110010111010110011101100100010111110110011101101000100001001001111010000100001111010000110000000011000000110000010100010100001011110100001101001000010010000100111001001010010010100100101001001001010011000100110101001001010010010100100101000111010001100100010101000110010001110100010101000100010001010100011001001000010010100100101001001011010010110100101101001110010100000101001001010100010101110101101001011011010111000101101101011101010110110101100101010110010101000101000001001111010011010100101001001001010001110100011001000100010000110100001001000010010001010100001001000101010001100100011101001001010010010100101101001110010011000100101101001010010011000100111101001011010010010011111100101011000101000000110000000111000001110000100100011011010101111001010110010101011110010110010001100000011001000101110001011011010111110110011001011111011000100101111001001111010100010100100000111011,
	960'b001010010011100001000010010000110100111101010110010101010110010101101100011000000101101001100101011000010101110101100011011001000110100110010100101001111000010101001000000110010000011100000011000001000000011100000100001011001011110001100111000001000000011100001101100100101010010000010110000010000000101000001001000001110001010110101000100100100000110100001001000010100000101000001011000010010001011010100111100100100000111100001010000010100000101000001001000010010000111010010101101000100001010100001001000010110000101100001010000001110000011110000100101100110010001000000111000010100000101000001001000010010000010101101010101111100010110000000110000010000000011000000110000010111001001010100011000101010000011000000010010100111100001000111101000000010000011000000101000001010000011100001101001010100101110110010010100110000111110001110011011010110110011101011011011000010110010001011000011001100110000101011100011010010110011101010100010001110100011000111111,
	960'b001011110011010000111011010001110100111001010011011000010110001101100110011001110110010001011010011000000110000001011011011000010110110001101101011110011001000010100011100101100111001101001001001010000001011000001011001000000111110001000111000001010000011000001011010111010110111100001101000001100000011000000110000001010000110101101001011000010000011100000111000010000000100000001000000001010000101101100111011000010000100000000111000001100000010000000101000001000000010101011100011011010000101000000010000000110000010000000100000000100000001101001101011110000001010000000100000001100000010100000110000001100000010101000000011111100010000100000100000001110000011000000110000010000101101101110000000011000000010100000101001101011000001000101100000001110001000000011110001101110101110110000101100111001001100001111101011011010110110001100110011001100110100001101010010111110101101001011100011000010110010001101010011000000101111001011100010100000100010000111110,
	960'b001100000011010100111010010010000100100001010010011001100110001001100100011010000110100101011100011000000110001001011111011001100111001101100011011001110110111001110100011110111000110010011100100111001001001110001000011101010110100101101001011010000110100101101000011001000110001101101011011010100110101001101010011010110110011101100101011001000110100101100111011011000110100101101001011010010110011101100011011001000110011101101001011010000110100101101001011010010110100001100100011001000110100001100110011010000110100001101001011010010110100101100110011000010110010101101000011001110110010101100111011010100110011101100100011001000110011101101010011010100110100001101000011010110110010101100101011010010110011101101000011001100110011001101101011111011000110110011000100111111001110110000111011100110110100001100010010111100110101001100101011001110110100001101010011000000101111001011100011000000110010101101011011001000101111101011010010011110100001100111110,
	960'b001010000011010101000000010000110100101101010001010110010110011101101000011001000101111001011111011000100110010001100101010111110110001101101100011010010110011001011101011000110110011101101100011100110111100010000110100101011001100010010010100100001001001010010000100100011001000110001111100101001001110010011001100100001001001010010110100100101001010110010011100100001001101010011010100101001000111110010000100101011001001010010101100100001001001010011011100110111001001110001110100101001001001010001110100100101001000010010010100110111001100110010001100100001001010010001110100100101001000110001101100100111001100110011001100100001001010110001101100010111001000110010001100100011001101110011001100011111001001010010010100100001001010110010011100001111000100110000110011110000110010001100101011001110110000001100100011000000101101001101000011010100110100101011100011000100110001001011101011000110110000101011100011010110110010101010010010011000100100101000001,
	960'b001010100011011100111101010000010100100101011001010110110110000101101001011000010110010101100111010111100110001001100101011010000110000001101100011010110101110101100101011001100110000101100000011001100110010001011111011010100110100001100101011011000110100001100011011001010110011101100101011001010110111101100110011001010110101001100110011001110110101001101100011001000110011101101111010111110110011101101011011000110110010001101010011011000110001001101011011100000110001101100110011010010110001001100010011000110110100101100100011011010110101101100001011010100110011001100010010111110110001101100111011000110110111101100100011000000110001001100000011000000110000101101001011000110110100001100111011001110110110001100101011001100110011001101010011010000110001101101100010111110110010001101000011000100110001101100000011010000110000101011111011001110110000101100101011001110110000101100011011000010110011001100010011000010101110001010000010100110100011001000000,
	960'b001011010011001000111101010011000100101001010010010111110101111001011111011000010110011101011110011001100110110001100001011000110110010101100001011000110110001101100111010111010110101001101001010111100110010101100110011000110110000001100111011000110101110101101010011001110101111101100110011000000110001101011101011001110110000001100011011011100110010001100010011001100101111001100010010111100110100101011111011001010110101101011110011000100110010001011101010111110101111001100111010110110110011101101100010111000110001001100101010111110101111101100010011000000101101101101010011001110101100101100110011000100110000001010111011000100101110001100010011000110101011001100010011000100101111101100000011001010101111001011111011011010110011101011101011001100110001101100001011000000110011001011011011001000111000101011111010111010110011101100010011000010110000101100110010110110110011001101111011000000110000101100100010111100101100101011000010100000100001001000011,
	960'b001010100011001100111100010010100100110001010100010111000101110101011100011010000110001101100100011001100110101001100011011000000110011101011101010110100110001101011011010111100110101001101010011000000110000101100100010111000101111001100100010111000101111001100111011001100110000101100001011001010101110101100100011001000101111101100100011011000110010101100000011000110110000101011011011001010110000101011101011001010110101001100001010111100110000001011011010110100110001101100000011000010110011101101010011000100110000101100101010111000101111001100101010111110110001001100101011000110101111101011110011001000101100001011000011000100110000101011101011000000110000101100001011000100101110001100000011000110110010101101100011010000110011001100011011000100110000101011000011000000101111001011110011001000110100101100101011000110110000101100001010111000110000001100001011000100110010001101010011001110110000101011110010110110101011001010111010011010100101101000001,
	960'b001010100011101001000011010001000101011101011010010101100101100101100011010111010110000101101111011010100110001101101101011001110101110101011011010111100101110001100000011011010110010101100100011011110110001001011010010111110110001101011101011010000111000001100100011011000110111101011110010110110110011001011110010111000110011101101110011000100111000001101010010111000101110001100010010111000101111001101011011000110110001001110001011001010101100001011010011001000101111101100010011011110110011101100110011011110110010001011010010111100110001001011011011000100111000101100011011000110110110101011111010110000101111101011011010110010110011001100000011001000110101001100001010110110110001001100100010110110110011101101110011000110110100101101110011000110101101001011110010111100101110001100100011010100110000001101011011010110101110101011010011001000110000101011111011011000110101001100111011100000110011001011010010111000101101101010011010011100100111101000011,
	960'b001010100011010100111101010010110100111001010010010101010101100101011011011001010110000001011111011001000110100101100011011000010110001001011001010110110110001101011101011000000110100001100111010111100110000001100101010111010101110001100100011000010110001001100111011001010101111101011111011000010101110001100100011000110101111101100011011001110110000101100000011001000110000101011011011001000110000101011011011000110110010001100000010111010110001001011101010111100110001001100010010111110110000101100111010111110101101101100010010111010101110001100010010111000101111101101001011000110101100101011001010111010101011001011011011000100101101001100001011000110101110001011100011000000101110001011110011001000101111001100000011011010110010001011110011001010101110101011001010111100110000001011010011000010110110001100010010111110110010101100001010111100110000101100100010111100110001101101001010111110101110001100010010110010101010101010111010011110100011101000100,
	960'b001011000011010000111011010010110100101001001111010110100101010101010111010110100110010001011011011001000110101001011100011000010101110001011000010111000101110101011111010110000110011101100111010110000110001001100000011000010101110001100011011000110101110001100101011000000101100001100011010111000110000001011010011001010101110001011110011010100101100101011110011001010101100101011111010110110110010001010111011000000110010101010101010111100101111101011000010111010101101001100101010110010101110101100100010101100101111101011111010110110101101001011100011000010101011101101000011000000101011001100000010101100101110001010011010111100101100101011101010111100101100001100001010110100101101101010101011000110110001001011010011001110101111001011110011000010101011101011110010101100110001001011111010110100110011001011010011000010110010101011101011001000101101101100110010111110110000001100110010110100101111101011110010101110101011001010011010100010100001101000000,
	960'b001010000011010100111100010000010100100101010011010100100101110001100001010110010101101001011110010101110101100101011110010111100101100001100000010111100101010101011101010111110101011101010111011000000101110101010110011001110110010001011001011000000101110101011001010101100110000001011011010110000110010101011100010110000101111001011001010110000101101101100001010110100110001101100110010110010101101001100001010101110101010101011100011000000101010001100001011001010101100001011010010111010101011101010110010111010110001001010111011000000110000001010100010111010101101101010110010101100101101101010101010101100110000101011000010100110101110101010111010101110101111101011001010101110110010001100000010100110101101101011010010101000101111001100001010101110101110101100010010111100101010101011100010111000101010101011010010111010101010101100001011010100101111101011000011000010101110001011000010111100101111001010101011000000101110101001011010011000100010100111000,
	960'b001001000010111100111001001111110100100101001100010100100101101101011111010110110101010001011000010101000101001101010100010100110101100001011101010111010101011101010000010101100101010101010100010101100101001101011010011000010110000101010111010100010101011001010110010101100101001101010011010110010110000001011110010101000101001101010111010100110101100101010000010101110101111101011110010111000101001001010010010101100101001001011010010011110101100001011110010111100101110101010010010100110101100001010011010101000101001001010110010111010101110101011000010011110101001101001111010100100101000001010010010110000101101001011000010101000101011001010101010101010101010101010111010110110101111001011011010110000101010001010100010100100101010101010010010110010101101001011011010110100101100101001110010101100101001101010100010100010101101001011100010111110101111001011000010100110101010101010110010101010101000101011010010110110101011101001111010001100011111100110100,
	960'b001001010010110100110011001111010100000001001100010101000101000001010011010101100101101001010010010011010100110101001101010101110101101101010000010100100101011001011001010100010100110101001100010100000101110001011000010100100101001001011011010101010100111101010000010011100101001101011101010101110101010001010110010111000101011001001101010011010100111001010100010111000101011001010100010101010101101101010010010011110100110101001101010101100101011101010010010100100101010001011001010011100101000001010000010011100101100001011011010100100101000101011000010101110100110101001100010010010100111001011001010100110100111001010010010101110101000001001111010011100101000001011100010101110101001001010010010110010101100001001110010011110100110001010011010111000101001001010000010101000101101001010101010011100101000001001100010101100101101101010001010100110101011001011100010100010100111101010000010011110101100001011011010100100100110101001111010010110011101100110000,
	960'b001000010010011000101111001101110011101101000011010010100100101001001100010011010100110101001000010010010100100101001000010010100100111001001011010010110100111001001011010010000100100001001000010001100100101101001100010011000100110001010000010010010100100101000110010010000100100001001101010011100100111001001101010011110100011101001000010010100100110001001001010100100101000001001111010011110100110101001000010001110100101001001010010010010100111101001110010011110100110001001001010001100100011101000100010010000100011001001111010011000100101001001111010010110100011001001000010001000100001101001001010011000100101001001010010011100100100101000110010001110100011001001010010010110100111001001101010010110100100001001001010001100100100101000111010010110100110101001011010011000100110001000110010001110100100001001001010001100100110001001111010011100100110101001010010001110100101001001000010010010100011001001101010011010100101101000011001110100011011100101111,
	960'b000111010010010100101100001100000011101000111010001110010100010101001000010001000011111001000101010000110100000101000101010000000100000001001011010010000100000101000011010001010100000001000010010001110011111101000001010011000100100000111111010001000100011000111110010001000100001100111101010001000100111101001000001111100100010101000101010000000100101001000100010000010100101001001011010001000100000001000100010000110100001101000101001111100100000001001010010010100100000100111111010001010100010001000000010001100100000000111110010011000100110001000001010000100100010100111110010000000100010000111101010000000100101101001000001111010100001101000000010000100100011001000000010000100100100101001001001111110100010001000011001111100100001001000100001111110100011101001011010001110100000101000111010001010011111001000111010001100011111001001001010010100100000100111110010010000100001100111111010001100100001000111111010001100100010100111010001101100011010000101000,
};

always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = r_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		g_data = g_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		b_data = b_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule