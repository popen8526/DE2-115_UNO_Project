module red_zero(
    input [7:0] addr,
    output [239:0] data
);
parameter [0:149][239:0] picture = {
    240'b111111101111111011111011101100001000000101100110010100000101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100111001010110100111110101111110111111110,
    240'b111111011111100111110011111101111111110011111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110011111001111101001111010111111100,
    240'b111111001111010011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111010111110101,
    240'b110111101111100111111111111111101111110111111001111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111110111111110111111111111110111110001,
    240'b100101011111111111111111111110101111100111111010111111001111101011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111010111111101111111111110111,
    240'b110101111111111111111101111110011111101011111110111111111111111011111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111101,
    240'b111110101111111111111101111110011111111011111100111110101111110111111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111111011111100111110011111110011111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111111011111100111110011111110011111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111111011111100111110011111110011111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111111011111100111110011111110011111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111111011111110111111011111111011111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111011111111011111110111111100111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111101011111110111111101111111011111010111110011111100111111001111110011111100111111001111110101111101011111101111111101111111011111111111111111111111111111111111111101111101011111001111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110011111101011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111010111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111101011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111010111111101111111111111111111111101111110011111100111111001111110011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111101111111111111111111111101111110101111100111111001111110011111100111111001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111110111111111111111111111111011111001111110011111100111111010111110111111100111111001111110011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111001111111001111111111111111111111111111110011111001111110101111110011111110111111111111110111111010111110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111001111111101111111111111111111111111111101011111001111110101111111111111111111111111111111111111100111110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111,
    240'b111110001111111111111101111110011111100111111100111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111101011111110111111111111111111111111111111111111111111111110111111101111111111111111,
    240'b111110001111111111111101111110011111100111111110111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111100111111101111111111111111111111111111111111111111111111100111111011111111111111111,
    240'b111110001111111111111101111110011111101011111111111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111100111111101111111111111111111111111111111111111111111111100111111011111111111111111,
    240'b111110001111111111111101111110011111111011111111111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111100111111101111111111111111111111111111111111111111011111001111111011111111111111111,
    240'b111110001111111111111101111110101111111111111111111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111100111111101111111111111111111111111111111111111110011111001111111011111111111111111,
    240'b111110001111111111111101111111001111111111111111111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111100111111101111111111111111111111111111111111111101011111001111111011111111111111111,
    240'b111110001111111111111101111111011111111111111111111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111101111110011111101011111111111111111111111111111111111111001111100111111001111111011111111111111111,
    240'b111110001111111111111110111111101111111111111111111111111111111111111111111111111111101011111001111110101111111111111111111111111111111111111100111110011111101011111111111111111111111111111111111110111111100111111001111111011111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111110011111101111111101111111111111110011111001111110011111101111111111111111111111111111111011111110011111100111111001111111011111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111111011111010111110011111100111111001111110101111100111111001111110101111111011111111111111111111110011111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111111100111111001111110011111100111111010111111101111111111111111111111111111101111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101111111011111110111111110111111111111111111111101111110111111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110011111100111111001111110011111100111111001111110011111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111111011111111111111111111111111111111111111111111111111111111111111111111111111111110111110111111101011111001111110011111100111111001111110011111100111111010111110101111100111111001111111011111111111111111,
    240'b111110001111111111111101111110011111101011111101111111101111111111111111111111111111110111111101111111011111110011111001111110011111100111111001111110011111100111111001111110011111110111111111111111111111101111111001111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110101111101111111011111110111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111001111111111111100111111011111111011111001111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111101111110111111001111110011111111011111100111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111101111110011111001111110011111111011111101111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111101111110011111001111110011111111011111101111111011111111111111111,
    240'b111110001111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111101111110011111001111110011111111011111101111111011111111111111111,
    240'b111110011111111111111101111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111100111111011111111011111001111111011111111111111111,
    240'b110000011111111111111110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111110111111111111111011111101111111001111111011111111111111011,
    240'b100111001111111111111111111110111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111010111110101111100111111011111111111111111111110100,
    240'b111100101111100111111111111111111111111011111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111111011111111111111111111101111110011,
    240'b111111101111011011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111111011,
    240'b111111011111110111010001110010001111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111001111100001111011111111101,
    240'b111111101111111011111011101100001000001001100110010100000101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100111001110110100111110101111110111111110,
    240'b111111011111100111110011111101111111110011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011111010111101001111010111111100,
    240'b111111001111010011111100111111111111111111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111111111111111101111010111110101,
    240'b110111101111100111111111111011011011101001110100011100110111011001111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011101111011011111101001111111111111110111110001,
    240'b100101011111111111101101100001110101100110000010101001100111111101011011010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101110010000010111010101111111111110111,
    240'b110101111111111111010100010111011000001011100111111110111110010001111111010111110110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011100110010101111111111111101,
    240'b111110101111111111010010011001101101111010111011011100101100001011011001011001010110000001100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011110110010001111111111111111,
    240'b111110001111111111010010011010111110110110100011010100101010101111101000011010010110000001100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011110110001111111111111111111,
    240'b111110001111111111010010011011011110110110100101010101011010110011101000011010010110000001100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011110110001111111111111111111,
    240'b111110001111111111010010011011011110110110100100010101011010110011101000011010010110000001100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011110110001111111111111111111,
    240'b111110001111111111010010011010101110101110100101010100011010110111100111011010000110000001100001011000010110000101100001011000010110000101100000011000000110000001011110010111000101110001011101011000000110000101011110110001111111111111111111,
    240'b111110001111111111010010011001001101111011100011101111011110010111011010011001000110000001100001011000010110000101100001010111100101111001100100011010010110100010010101101110111011101110101100011010100101111101011110110001111111111111111111,
    240'b111110001111111111010011010111011000101011100000111010101101111010000111010111110110000101100001011000010101111101011111011101101000011011010010111001011110011111110101111111111111111111111101111001001001000101011010110001111111111111111111,
    240'b111110001111111111010011010111110101111101100110011010000110011001100000011000010110000101100000010110110111001010100110111011011111110011111111111111111111111111111111111111111111111111111111111111111111000010000101110000111111111111111111,
    240'b111110001111111111010011010111110110000101100000011000000110000001100001011000010101111101100011101000011101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011110111011111111011111111,
    240'b111110001111111111010011010111110110000101100001011000010110000101100001010111010111101111010100111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111110111111111,
    240'b111110001111111111010011010111110110000101100001011000010110000101011101011101101101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111011111111,
    240'b111110001111111111010011010111110110000101100001011000010101111001110001110110011111111111111111111011111010100010011100100111011001111011000001111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111,
    240'b111110001111111111010011010111110110000101100001010111110110101011001111111111111111110111000110011110100101111001010111010101100101100101100101110000001111111111111111111111111111111111111111111111111111111111111111111110111111111011111111,
    240'b111110001111111111010011010111110110000101011111011001001100001011111111111111111110110101110000010110110101110001111110100100000110111001011100011010001100110111111111111111111111111111111111111111111111111111111111111100111111111011111111,
    240'b111110001111111111010011010111110110000101011111101011111111111111111111111111111011010001011111011001111010101111101000111111111100100001101000010110111000100011111101111111111111111111111111111111111111111111111100111011101111111011111111,
    240'b111110001111111111010011010111110101111101101111111001111111111111111111111111111000100001011010011101011111011111111111111111111111111110110110010110101000010011111011111111111111111111111111111111111111111111111011111100001111111011111111,
    240'b111110001111111111010011010111110101101010101110111111101111111111111111111111001000100101011011011110111111011111111111111111111111111111001100010110110111100011101001111111111111111111111111111111111111111111100111111000011111111011111111,
    240'b111110001111111111010011010111010111001011011111111111111111111111111111111110111000100001011011011111111111100011111111111111111111111111001010010111100101111010111110111111111111111111111111111111111111111110111100110000111111111111111111,
    240'b111110001111111111010011010111001001011011111111111111111111111111111111111110111000100001011011011111111111100011111111111111111111111111001010010111100101111110111111111111111111111111111111111111111111111010101101110000101111111111111111,
    240'b111110001111111111010010011000111101110011111111111111111111111111111111111110111000100001011011011111111111100011111111111111111111111111001010010111100101111110111111111111111111111111111111111111111110111001101110110001011111111111111111,
    240'b111110001111111111010000100011001111010111111111111111111111111111111111111110111000100001011011011111111111100011111111111111111111111111001010010111100101111110111110111111111111111111111111111111111011101101011110110001111111111111111111,
    240'b111110001111111111001110101110011111111111111111111111111111111111111111111110111000100001011011011111111111100011111111111111111111111111001010010111100110000111000011111111111111111111111111111110011000001101011010110001111111111111111111,
    240'b111110001111111111001111101111101111111111111111111111111111111111111111111111011000101001011011011110101111011111111111111111111111111111001100010110100111111011110011111111111111111111111111110000100110000101011101110001111111111111111111,
    240'b111110001111111111100010110110011111111111111111111111111111111111111111111111111000101001011010011100111111001011111111111111111111101110100010010110101000010011111011111111111111111111110011100011000101110101011110110001111111111111111111,
    240'b111110001111111111111000111101101111111111111111111111111111111111111111111111111100100001100010011001001000101111010011111100111010111101100001010110111001000111111110111111111111101110011111010111010110000101011110110001111111111111111111,
    240'b111110001111111111111010111110001111111111111111111111111111111111111111111111111111000101111101010110100101110001101011011100100110010001011100011101111110000111111111111111111011111001100000011000000110000101011110110001111111111111111111,
    240'b111110001111111111111110111111101111111111111111111111111111111111111111111111111111111111011100100101100110001001011010010110100101101101110010110110001111111111111111111011101000011101011101011000010110000101011110110001111111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100101110111101101111011100010011011101111111111111111111001000100000100101111101100001011000010110000101011110110001111111111111111111,
    240'b111110001111111111111101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001101010010111000110000101100001011000010110000101011110110001111111111111111111,
    240'b111110001111111111101001111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101110100110111101011110011000010110000101100001011000010110000101011110110001111111111111111111,
    240'b111110001111111111001110101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110110010011010111000110000001100001011000010101111101011110010111100110000001011110110001111111111111111111,
    240'b111110001111111111010001011100011101011111111111111111111111111111111111111111111111111111111111111111111111011111011000100010010111010101100000011000000110000101100001010111110110110001111111011111000110010001011101110001111111111111111111,
    240'b111110001111111111010011010111000111100010111111110101011111110111111101111111111101011111000101110000011001101101100100010111110101111001100001011000010110000101011111011010011100100111111100111110011010100101011110110001111111111111111111,
    240'b111110001111111111010011010111110101111101011100011011001001011110010111100110010110111001011101010111000101110101100000011000010110000101100001011000010110000001100000101110011111100110101000110000111110110001101010110001011111111111111111,
    240'b111110001111111111010011010111110110000101100001010111110101110001011100010110110101111101100001011000010110000101100001011000010110000101100001011000010110000001100011111000101100001101011101011010111110000110100110110000101111111111111111,
    240'b111110001111111111010011010111110110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000001100011111000011011100101011100011000101101111010110110110000011111111111111111,
    240'b111110001111111111010011010111110110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000001100011111000101011100101011100011000101101111010110101110000011111111111111111,
    240'b111110001111111111010011010111110110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000001100010110101111100000001011100011010011110000110101011110000011111111111111111,
    240'b111110011111111111010011011000000110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011101100011011111100010100101110000111110110101101011110001111111111111111111,
    240'b110000011111111111010110011000010101111001100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111011010111100101111111111110110111001011101011111110011101111111111111011,
    240'b100111001111111111110110100111110110100001011110010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111000110101110000001011011110110001010011000111101001111111111110100,
    240'b111100101111100111111111111110111101011010011001100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001100110010111100110001101010011111000111111111111101111110011,
    240'b111111101111011011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111111011,
    240'b111111011111110111010001110010001111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111001111100001111011111111101,
    240'b111111101111111011111011101100111000010101101000010100000101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100111010010110101111110101111110111111110,
    240'b111111011111100111110011111101111111110011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011111010111101001111010111111100,
    240'b111111001111010011111100111111111111111111110110111101101111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101101111111111111111111111101111010111110101,
    240'b110111101111100111111111111011011011011101101110011011010111000001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011100101011010111101001111111111111110111110001,
    240'b100101011111111111101100100000100101001101111101101000100111101001010100010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101010101111100111010011111111111110111,
    240'b110101111111111111010010010101100111110111100110111110111110001101111001010101110101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100101010100110010001111111111111101,
    240'b111110101111111111001111010111111101110110111000011010111011111111011000010111100101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111001111011001011110110010011111010010111010011111101000011000110101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111001111011001111110110010100000010011101010100111100111011000110101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111001111011001111110110010011111010011101010100111100111011000110101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111001111011001001110101110100000010010011010100111100111011000100101100101011010010110100101101001011010010110100101101001011001010110010101100101010111010101010101010101010101010110010101101001010110110001011111111111111111,
    240'b111110001111111111010000010111011101110111100010101110101110010011011000010111010101100101011010010110100101101001011010010101110101011101011110011000100110001010010000101110011011100010101000011001000101100101010110110001011111111111111111,
    240'b111110001111111111010001010101101000010111011111111010011101110110000001010110000101101001011010010110100101011101011000011100001000000111010001111001001110011011110101111111111111111111111101111001001000110101010011110001011111111111111111,
    240'b111110001111111111010001010110000101100001100000011000100101111101011001010110100101101001011001010101000110110010100011111011001111110011111111111111111111111111111111111111111111111111111111111111111110111110000000110000011111111111111111,
    240'b111110001111111111010001010110000101101001011001010110010101100101011010010110100101100001011100100111011101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110111001111111011111111,
    240'b111110001111111111010001010110000101101001011010010110100101101001011010010101010111011011010001111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111110111111111,
    240'b111110001111111111010001010110000101101001011010010110100101101001010110011100001101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111011111111,
    240'b111110001111111111010001010110000101101001011010010110100101011101101010110101111111111111111111111011101010010110011001100110011001101010111110111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111,
    240'b111110001111111111010001010110000101101001011010010110000110001111001100111111111111110111000100011101010101011101010000010011110101001001011110101111101111111111111111111111111111111111111111111111111111111111111111111110111111111011111111,
    240'b111110001111111111010001010110000101101001011000010111101011111111111111111111111110110001101010010101010101010101111001100010110110011101010101011000101100101111111111111111111111111111111111111111111111111111111111111100111111111011111111,
    240'b111110001111111111010001010110000101101001011000101010111111111011111111111111111011000101011001011000011010011111101000111111111100011001100010010100111000010011111101111111111111111111111111111111111111111111111100111011101111111011111111,
    240'b111110001111111111010001010110000101100001101000111001101111111111111111111111111000010001010011011100001111011111111111111111111111111110110010010100100111111011111011111111111111111111111111111111111111111111111011111100001111111011111111,
    240'b111110001111111111010001010110000101001110101010111111101111111111111111111110111000010001010011011101101111011111111111111111111111111111001010010101000111001011101000111111111111111111111111111111111111111111100110111000001111111011111111,
    240'b111110001111111111010001010101100110110011011110111111111111111111111111111110111000001101010011011110101111100011111111111111111111111111001000010110000101011110111011111111111111111111111111111111111111111110111001110000001111111111111111,
    240'b111110001111111111010001010101011001000111111111111111111111111111111111111110111000001101010011011110101111100011111111111111111111111111001000010110000101100010111100111111111111111111111111111111111111111010101010110000001111111111111111,
    240'b111110001111111111001111010111001101101111111111111111111111111111111111111110111000001101010011011110101111100011111111111111111111111111001000010110000101100010111100111111111111111111111111111111111110110101101000110000111111111111111111,
    240'b111110001111111111001101100010001111010111111111111111111111111111111111111110111000001101010011011110101111100011111111111111111111111111001000010110000101100010111011111111111111111111111111111111111011100001011000110001011111111111111111,
    240'b111110001111111111001100101101101111111111111111111111111111111111111111111110111000001101010011011110101111100011111111111111111111111111001000010110000101101011000000111111111111111111111111111110000111110101010010110001011111111111111111,
    240'b111110001111111111001101101110111111111111111111111111111111111111111111111111001000010101010011011101011111011111111111111111111111111111001011010100110111100011110011111111111111111111111111101111110101101001010110110001011111111111111111,
    240'b111110001111111111100000110101111111111111111111111111111111111111111111111111111000011001010011011011101111001011111111111111111111101110011101010100100111111111111011111111111111111111110011100001100101011001010110110001011111111111111111,
    240'b111110001111111111111000111101101111111111111111111111111111111111111111111111111100011001011011010111011000011011010010111100111010101101011010010101001000110111111110111111111111101110011100010101100101101001010110110001011111111111111111,
    240'b111110001111111111111010111110001111111111111111111111111111111111111111111111111111000101111000010100110101010101100100011011010101110101010101011100011110000011111111111111111011101101011001010110010101101001010110110001011111111111111111,
    240'b111110001111111111111110111111101111111111111111111111111111111111111111111111111111111111011011100100100101101101010011010100110101010001101100110101101111111111111111111011011000001001010110010110100101101001010110110001011111111111111111,
    240'b111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100100110111011101110111100000111011100111111111111111111000111011111100101011101011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111111101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101001100101010101010101101001011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111100111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000101101110110100101010111010110100101101001011010010110100101101001010110110001011111111111111111,
    240'b111110001111111111001011101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110010001111010101010101100101011010010110100101100001010111010101110101100101010110110001011111111111111111,
    240'b111110001111111111001111011010101101011011111111111111111111111111111111111111111111111111111111111111111111011111010111100001000111000001011001010110010101101001011010010110000110010101111010011101110101110101010101110001011111111111111111,
    240'b111110001111111111010001010101000111001010111100110100111111111011111110111111111101010111000011101111101001011101011101010110000101011101011010010110100101101001011000011000101100011111111100111110011010010101010111110001011111111111111111,
    240'b111110001111111111010001010110000101100001010101011001101001001110010011100101010110100001010110010101010101011001011001010110100101101001011010010110100101100101011001101101101111101010100100110000011110101101100100110000111111111111111111,
    240'b111110001111111111010001010110000101101001011010010110000101010001010100010101000101100001011010010110100101101001011010010110100101101001011010010110100101100101011100111000011100000101010110011001011110000010100011110000001111111111111111,
    240'b111110001111111111010001010110000101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100101011100111000001011010001010101010111001101110010110010101111111111111111111111,
    240'b111110001111111111010001010110000101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100101011100111000101011010101010101010111001101110010110001101111111111111111111111,
    240'b111110001111111111010001010110000101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100101011011110101101011110101010101011001001101111110100111101111111111111111111111,
    240'b111110011111111111010010010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010110100010001111100010100001110000001110110101100101110001001111111111111111,
    240'b110000011111111111010101010110100101011101011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011000011001011100100011111111110110011001001101010111110010111111111111111011,
    240'b100111001111111111110110100110110110000101010111010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010101010110010001111100011010010101101110010100111101001111111111110100,
    240'b111100101111100111111111111110111101010110010110100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100110001001011010010011100101001101001111111000111111111111101111110011,
    240'b111111101111011011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111111011,
    240'b111111011111110111010001110010001111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111001111100001111011111111101,
    };
    assign data = picture[addr];
endmodule