module blue_eight(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111111111111110111100100101000101010001011000000110000111100001111000011110000111100001111000010110000101100001011000010110000101100001111000011110000111100001111000011110000101100001011000011101111011001110110110101111110001111111111111111,
	240'b111111111111100010111111110001001110000111100100111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001101111111000010110100101111111011111111,
	240'b111111111100101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011011101011111111110,
	240'b110100011100110111111111111110101100010010100100101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010011110101001011100111011111110111111011100011011001101,
	240'b100110001110110011111111101010100101001101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110110001001110100010101000101011111000001111111111101111010011000,
	240'b101001001111100011110011011010100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011011101101111111110100101100110101000001111111111111011110100110100110,
	240'b101101011111110011101001011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111101001101110000110100011111011110110011101110000111110011110111010110111,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111100101101110110011001001111001100101111101110000111110011110111110111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101011101111100111101011111100000111010101101111111110011110111110111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010111001100101100000110100101011011101101111111110011110111110111000,
	240'b101101101111110011101001011000010101001101010100010100000101000001010000010100000101000001010010010101000101010101010101010101010101010101010101010101010101001001101111111011110111110001001000101111101100010001110000111110001110111110111000,
	240'b101101101111110011101001011000010101000001011101100000111001101110011010100100000111111001101001010101100101000001010010010101010101010101010101010101010101010001011001110100101101111010110101111101011001001101101110111110011110111110111000,
	240'b101101101111110011101001010111010111000111010010111111001111111111111111111111111111101011101011110011011010000101110000010100110101001001010101010101010101010101010010011100001100101111100010101010000101010101110010111110011110111110111000,
	240'b101101101111110011100111011100101101111011111111111111111111111111111111111111111111111111111111111111111111111111110000101110000111000001010001010101000101010101010101010100100101011101011110010100110101000101110011111110011110111110111000,
	240'b101101101111110011100101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110011111010110010101001001010101010101010101010001010011010101010101001001110011111110011110111110111000,
	240'b101101101111101011110001111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110110010001010001010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111100111111010111111001111111111111111111111111111111111111111111111111111111111111111111111111111110111101110111100001111111111111111111111111101011001101100010100010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111100111111010111111011111111111111111111111111111111111111111111111111111111111111111111001011000110101100100011001111001101111110000111111111111111111011010011010100101000101010101010101010101001001110011111110011110111110111000,
	240'b101101101111100111111001111110011111111111111111111111111111111111111111111111111111111111110001011110110100111001001110010011100100111010001111111110101111111111111111110100000101111001010011010101010101001001110011111110011110111110111000,
	240'b101101101111101011110100111011111111111111111111111111111111111111111111111111111111111110111001010100000101010101111110011101100101001101010110110100101111111111111111111111111011001101010011010101000101001001110011111110011110111110111000,
	240'b101101101111101111101100110111101111111111111111111111111111111111111111111111111111111110010101010011000111011111110111111010000110010101001101101100011111111111111111111111111111100110001000010100000101001001110011111110011110111110111000,
	240'b101101101111101111100101110001111111111111111111111111111111111111111111111111111111111110010101010011000111011111111000111010010110010101001110101100001111111111111111111111111111111111011011010111100101000001110011111110011110111110111000,
	240'b101101101111110011100100101001011111111111111111111111111111111111111111111111111111111110111101010100110101010101111110011101100101001101011010110101011111111111111111111111111111111111111111100110110100110001110011111110011110111110111000,
	240'b101101101111110011100101100000101111011011111111111111111111111111111111111111111111111111010011010110110101001101001111010100000101001001100111111001111111111111111111111111111111111111111111110111010101101001110001111110011110111110111000,
	240'b101101101111110011101000011001101101011111111111111111111111111111111111111111111111000101111001010100010101001101011111010111100101001001010001100011011111101011111111111111111111111111111111111111011000011001101110111110011110111110111000,
	240'b101101101111110011101001010111001010010011111111111111111111111111111111111111111011010101010000010101001001101011100000110111001000101001010001010101101100111011111111111111111111111111111111111111111011101101110000111110011110111110111000,
	240'b101101101111110011101001010111010110110011110001111111111111111111111111111111011000011101001100011111011111100111111111111111111110110001101001010011001010000111111111111111111111111111111111111111111110010010000001111101111110111110111000,
	240'b101101101111110011101001011000000101000110110111111111111111111111111111111110000111011001001100101000111111111111111111111111111111111110001000010010111000111011111111111111111111111111111111111111111111100110011100111101011110111110111000,
	240'b101101101111110011101001011000010101000001101110111011111111111111111111111110110111110101001100100101011111111111111111111111111111110001111100010010111001011011111111111111111111111111111111111111111111111110111101111100111110111110111000,
	240'b101101101111110011101001011000010101001101010001101000101111111111111111111111111001110001001101011000101101010011111111111111111100000001011000010011111011011011111111111111111111111111111111111111111111111111010110111101001110111010111000,
	240'b101101101111110011101001011000010101001101010011010110111101000111111111111111111101011101011011010100000110010110010111100100000101111001001111011010011110100111111111111111111111111111111111111111111111111111100101111110011110111010111000,
	240'b101101101111110011101001011000010101001101010101010100010111000011100111111111111111111010101101010101010100111001001110010011100100111001011100110000111111111111111111111111111111111111111111111111111111111111101111111111001110111010111000,
	240'b101101101111110011101001011000010101001101010101010101010101000010000000111011101111111111111101101111010111011001100001011000100111111011001100111111111111111111111111111111111111111111111111111111111111111111110100111111011110111010111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010000100001001110110011111111111111111111011011100011111001101111101011111111111111111111111111111111111111111111111111111111111111111111111111110011111111011110111010111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010100010111011111011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111110001110111010111000,
	240'b101101101111110011101001011000010101001101010101010101000101010101010101010101010101000101100101101110101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101111101001110111110111000,
	240'b101101101111110011101001011000010101001001010010010110100101001101010011010101010101010101010010010101011000001111001100111110001111111111111111111111111111111111111111111111111111111111111111111111111100111001111011111101111110111110111000,
	240'b101101101111110011101001010111110101101110101101110101111011001001100000010100110101010101010101010101000101000001011000011111101011011011011111111101101111111111111111111111111111111111111110110011110110011101101111111110011110111110111000,
	240'b101101101111110011101001010111011010011111110010110000001111000010110011010100110101010101010101010101010101010101010100010100010101001001011111011101111000110110100001101010111010100010001000010111000100111101110011111110011110111110111000,
	240'b101101101111110011101000011000111101111010100110010001111001101011100111010111000101010001010101010101010101010101010101010101010101010101010011010100010101000001010001010100010101000101010001010101000101001001110011111110011110111110111000,
	240'b101101101111110011101000011000101101011010110101010101101010110011100000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111110011101001010111011001000111110110110111111111011110011100010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111110011101001010111010111000111101111110100111111000101111010010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111110011101001010110111000000011101110100100111110101110001100010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110010111110011110111110111000,
	240'b101001101111100111110001011001100101110011010001111101111101100001100100010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001111100111111001110100110101001,
	240'b100101101110110111111110101000100100111101011111100000010110001001001110010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110101010110111010111111111101111110010110,
	240'b110010111101000011111111111101111011011110010101100100111001011010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001100001111111101111111101100011111000111,
	240'b111111011100011011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101001011111100,
	240'b111101001111000011000101110011111110001111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110001011000111110001011111001011110100,
	240'b111011101111010111110100101001111001000110101111101100111011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110011101011001000110010101011111011001111000011101111,
	240'b111111111111110111100100101000101010001011000000110000111100001111000011110000111100001111000010110000101100001011000010110000101100001111000011110000111100001111000011110000101100001011000011101111011001110110110101111110001111111111111111,
	240'b111111111111100010111111110001001110000111100100111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001101111111000010110100101111111011111111,
	240'b111111111100101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011011101011111111110,
	240'b110100011100110111111111111110101100010010100100101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010011110101001011100111011111110111111011100011011001101,
	240'b100110001110110011111111101010100101001101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110110001001110100010101000101011111000001111111111101111010011000,
	240'b101001001111100011110011011010100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011011101101111111110100101100110101000001111111111111011110100110100110,
	240'b101101011111110011101001011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111101001101110000110100011111011110110011101110000111110011110111010110111,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111100101101110110011001001111001100101111101110000111110011110111110111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101011101111100111101011111100000111010101101111111110011110111110111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010111001100101100000110100101011011101101111111110011110111110111000,
	240'b101101101111110011101001011000010101001101010100010100000101000001010000010100000101000001010010010101000101010101010101010101010101010101010101010101010101001001101111111011110111110001001000101111101100010001110000111110001110111110111000,
	240'b101101101111110011101001011000010101000001011101100000111001101110011010100100000111111001101001010101100101000001010010010101010101010101010101010101010101010001011001110100101101111010110101111101011001001101101110111110011110111110111000,
	240'b101101101111110011101001010111010111000111010010111111001111111111111111111111111111101011101011110011011010000101110000010100110101001001010101010101010101010101010010011100001100101111100010101010000101010101110010111110011110111110111000,
	240'b101101101111110011100111011100101101111011111111111111111111111111111111111111111111111111111111111111111111111111110000101110000111000001010001010101000101010101010101010100100101011101011110010100110101000101110011111110011110111110111000,
	240'b101101101111110011100101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110011111010110010101001001010101010101010101010001010011010101010101001001110011111110011110111110111000,
	240'b101101101111101011110001111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110110010001010001010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111100111111010111111001111111111111111111111111111111111111111111111111111111111111111111111111111110111101110111100001111111111111111111111111101011001101100010100010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111100111111010111111011111111111111111111111111111111111111111111111111111111111111111111001011000110101100100011001111001101111110000111111111111111111011010011010100101000101010101010101010101001001110011111110011110111110111000,
	240'b101101101111100111111001111110011111111111111111111111111111111111111111111111111111111111110001011110110100111001001110010011100100111010001111111110101111111111111111110100000101111001010011010101010101001001110011111110011110111110111000,
	240'b101101101111101011110100111011111111111111111111111111111111111111111111111111111111111110111001010100000101010101111110011101100101001101010110110100101111111111111111111111111011001101010011010101000101001001110011111110011110111110111000,
	240'b101101101111101111101100110111101111111111111111111111111111111111111111111111111111111110010101010011000111011111110111111010000110010101001101101100011111111111111111111111111111100110001000010100000101001001110011111110011110111110111000,
	240'b101101101111101111100101110001111111111111111111111111111111111111111111111111111111111110010101010011000111011111111000111010010110010101001110101100001111111111111111111111111111111111011011010111100101000001110011111110011110111110111000,
	240'b101101101111110011100100101001011111111111111111111111111111111111111111111111111111111110111101010100110101010101111110011101100101001101011010110101011111111111111111111111111111111111111111100110110100110001110011111110011110111110111000,
	240'b101101101111110011100101100000101111011011111111111111111111111111111111111111111111111111010011010110110101001101001111010100000101001001100111111001111111111111111111111111111111111111111111110111010101101001110001111110011110111110111000,
	240'b101101101111110011101000011001101101011111111111111111111111111111111111111111111111000101111001010100010101001101011111010111100101001001010001100011011111101011111111111111111111111111111111111111011000011001101110111110011110111110111000,
	240'b101101101111110011101001010111001010010011111111111111111111111111111111111111111011010101010000010101001001101011100000110111001000101001010001010101101100111011111111111111111111111111111111111111111011101101110000111110011110111110111000,
	240'b101101101111110011101001010111010110110011110001111111111111111111111111111111011000011101001100011111011111100111111111111111111110110001101001010011001010000111111111111111111111111111111111111111111110010010000001111101111110111110111000,
	240'b101101101111110011101001011000000101000110110111111111111111111111111111111110000111011001001100101000111111111111111111111111111111111110001000010010111000111011111111111111111111111111111111111111111111100110011100111101011110111110111000,
	240'b101101101111110011101001011000010101000001101110111011111111111111111111111110110111110101001100100101011111111111111111111111111111110001111100010010111001011011111111111111111111111111111111111111111111111110111101111100111110111110111000,
	240'b101101101111110011101001011000010101001101010001101000101111111111111111111111111001110001001101011000101101010011111111111111111100000001011000010011111011011011111111111111111111111111111111111111111111111111010110111101001110111010111000,
	240'b101101101111110011101001011000010101001101010011010110111101000111111111111111111101011101011011010100000110010110010111100100000101111001001111011010011110100111111111111111111111111111111111111111111111111111100101111110011110111010111000,
	240'b101101101111110011101001011000010101001101010101010100010111000011100111111111111111111010101101010101010100111001001110010011100100111001011100110000111111111111111111111111111111111111111111111111111111111111101111111111001110111010111000,
	240'b101101101111110011101001011000010101001101010101010101010101000010000000111011101111111111111101101111010111011001100001011000100111111011001100111111111111111111111111111111111111111111111111111111111111111111110100111111011110111010111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010000100001001110110011111111111111111111011011100011111001101111101011111111111111111111111111111111111111111111111111111111111111111111111111110011111111011110111010111000,
	240'b101101101111110011101001011000010101001101010101010101010101010101010101010100010111011111011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111110001110111010111000,
	240'b101101101111110011101001011000010101001101010101010101000101010101010101010101010101000101100101101110101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101111101001110111110111000,
	240'b101101101111110011101001011000010101001001010010010110100101001101010011010101010101010101010010010101011000001111001100111110001111111111111111111111111111111111111111111111111111111111111111111111111100111001111011111101111110111110111000,
	240'b101101101111110011101001010111110101101110101101110101111011001001100000010100110101010101010101010101000101000001011000011111101011011011011111111101101111111111111111111111111111111111111110110011110110011101101111111110011110111110111000,
	240'b101101101111110011101001010111011010011111110010110000001111000010110011010100110101010101010101010101010101010101010100010100010101001001011111011101111000110110100001101010111010100010001000010111000100111101110011111110011110111110111000,
	240'b101101101111110011101000011000111101111010100110010001111001101011100111010111000101010001010101010101010101010101010101010101010101010101010011010100010101000001010001010100010101000101010001010101000101001001110011111110011110111110111000,
	240'b101101101111110011101000011000101101011010110101010101101010110011100000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111110011101001010111011001000111110110110111111111011110011100010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111110011101001010111010111000111101111110100111111000101111010010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110011111110011110111110111000,
	240'b101101101111110011101001010110111000000011101110100100111110101110001100010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110010111110011110111110111000,
	240'b101001101111100111110001011001100101110011010001111101111101100001100100010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001111100111111001110100110101001,
	240'b100101101110110111111110101000100100111101011111100000010110001001001110010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110101010110111010111111111101111110010110,
	240'b110010111101000011111111111101111011011110010101100100111001011010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001100001111111101111111101100011111000111,
	240'b111111011100011011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101001011111100,
	240'b111101001111000011000101110011111110001111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110001011000111110001011111001011110100,
	240'b111011101111010111110100101001111001000110101111101100111011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110011101011001000110010101011111011001111000011101111,
	240'b111111111111110111100100101000101010001011000000110000111100001111000011110000111100001111000010110000101100001011000010110000101100001111000011110000111100001111000011110000101100001011000011101111011001110110110101111110001111111111111111,
	240'b111111111111100010111111110001001110000111100100111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001101111111000010110100101111111011111111,
	240'b111111111100101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011011101011111111110,
	240'b110100011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100011011001101,
	240'b100110001110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111010011000,
	240'b101001001111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010100110,
	240'b101101011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110110111,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101101101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110111000,
	240'b101001101111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010101001,
	240'b100101101110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110010110,
	240'b110010111101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011111000111,
	240'b111111011100011011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101001011111100,
	240'b111101001111000011000101110011111110001111100101111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001011110001011000111110001011111001011110100,
	240'b111011101111010111110100101001111001000110101111101100111011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110011101011001000110010101011111011001111000011101111,
};
assign data = picture[addr];
endmodule