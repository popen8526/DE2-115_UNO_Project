module red_four(
    input [7:0] addr,
    output [239:0] data
);
parameter [0:149][239:0] picture = {
    240'b111100101111101111010100101101011011011010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011010010110110110111011111001011101111,
    240'b111101001101000011001011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000101110011101101111110011,
    240'b110100101100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011100111100011,
    240'b101100011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100110100110,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010010111,
    240'b101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010101010,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
    240'b101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101011,
    240'b101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010011010,
    240'b101100011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010100001,
    240'b110010101101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011110011011100,
    240'b111100011100011111010111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110000001101000011110011,
    240'b111110001111010111000011101011111011110011000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011011110110010110101111111100011110110,
    240'b111100101111101111010100101101011011011010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011010010110110110111011111001011101111,
    240'b111101001101000011001011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000101110011101101111110011,
    240'b110100101100101011111111111111111111001111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100011101000111010101111101111111111111101001011100111100011,
    240'b101100011111010111111111110000100111010001100111011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001100110011010011000100011100101111111111101100110100110,
    240'b101101101111111111100010011000010100111101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010010010100101001100010010101010100000100110110001010111111011111001110010111,
    240'b101110101111111110111101010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100001001010111101000011001010101000001100110111011111111111010101010,
    240'b101111011111111110111000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110100011100011100111000100110101100101111010111111111110101110,
    240'b101111011111111110111000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000011100010010101111110110010101100101100011111010111111111110101110,
    240'b101111011111111110111000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111100011001110101001110010111001111000011001100000111010111111111110101110,
    240'b101111011111111110111000010100100101010101010101010101010101010001010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101101000001110111001111011110011111100011001100100111010101111111110101110,
    240'b101111011111111110111000010100100101010001010001010100010101010101010100010100010101000001010001010100110101010001010101010101010101010101010101010101010101001001100111111010011111111011110001111101111101101001101100111010011111111110101110,
    240'b101111001111111110111000010100010101010010000001101101011100010011000000101110001010000110000100011001100101010001010001010101000101010101010101010101010101010001011000101100001111011010010100100011010111111001100111111010111111111110101110,
    240'b101111001111111110110111010101001010110011110111111111111111111111111111111111111111111111111100111001111100000110000110010110010101000101010100010101010101010101010001011101101011001001010110010011110100111101100101111010111111111110101110,
    240'b101111001111111110110100100110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111011110011111000001001010100010100100101010101010101010101010101010001010101010101010101001101100101111010111111111110101110,
    240'b101111001111111111000101111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110110011000110101000101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111001111111111100001111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111001101010001010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111001111111111110000111111001111111111111111111111111111111111111111111111111111111111111111111110011101011011010010111010111111111111111111111111111110011001111010010100000101010101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111111101111111111001111111111111111111111111111111111111111111111111111111111111111111101110111111001001111100011011111110111111111111111111111111111100111011101010101000101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111111101010111110111111111111111111111111111111111111111111111111111111111111111111111111111011100001001111010111001101110011111111111111111111111111111111110111010110011001010010010101010101001101100101111010111111111110101110,
    240'b101111011111111111100001111110011111111111111111111111111111111111111111111111111111111111111111111111111110111101101100010011011001111011111111111111111111111111111111111111111100000101010111010101000101001101100101111010111111111110101110,
    240'b101111011111111111010100111101001111111111111111111111111111111111111111111111111111111111111111111111111111111110100110010011100110100011101010111111111111111111111111111111111111110110010101010100000101001101100101111010111111111110101110,
    240'b101111011111111111000111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011000000100111110110011111111111111111111111111111111111111111111100110011001100101000001100101111010111111111110101110,
    240'b101111001111111110111000110010011111111111111111111111111111111111111111111111111111111111101001100100101000101111011000100101000100110001110110111101011111111111111111111111111111111111111111101010010100111101100101111010111111111110101110,
    240'b101111001111111110110011101000101111111111111111111111111111111111111111111111111111111111011110010110010100110111000111110101100101011101010100110001101111111111111111111111111111111111111111111001110110001101100010111010111111111110101110,
    240'b101111001111111110110100011101101111100011111111111111111111111111111111111111111111111111011111010111100101001111000101111111010111111101001011100001101111110011111111111111111111111111111111111111111001010101100000111010111111111110101110,
    240'b101111001111111110110111010101111101011011111111111111111111111111111111111111111111111111011111010111100101001111000100111111111011111001010001010110111101100111111111111111111111111111111111111111111100101001100110111010101111111110101110,
    240'b101111001111111110111000010011011001101011111111111111111111111111111111111111111111111111100011010111100101001111000111111111111111011001110011010011001001100111111111111111111111111111111111111111111110111101111101111010001111111110101110,
    240'b101111001111111110111000010100000110010011100101111111111111111111111111111111111110101010111111010111000101001110101100110110111101110010010001010011110110010111101001111111111111111111111111111111111111110110011110111001101111111110101110,
    240'b101111011111111110111000010100100101000010011100111111111111111111111111111111111010000101010100010101010101010101011001010111000101110001011010010101000101011111011001111111111111111111111111111111111111111111000000111001101111111110101110,
    240'b101111011111111110111000010100100101001101011110110101011111111111111111111111111001100101001001010101010101010101010001010011100100111001001111010011110101001111011000111111111111111111111111111111111111111111011001111010111111111110101110,
    240'b101111011111111110111000010100100101010101010000011111001111010011111111111111111100100110001101010110010101010010000101101000001001111010011110100111101010000011101010111111111111111111111111111111111111111111101100111100011111111110101110,
    240'b101111011111111110111000010100100101010101010101010100011001110111111101111111111111111111100001010111100101001011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101011111111110101110,
    240'b101111011111111110111000010100100101010101010101010101000101010110110010111111111111111111011111010111010101001011000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111101101111111110101110,
    240'b101111001111111110111000010100100101010101010101010101010101001101011000101101111111111111110100110000101011111011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101111111111110101110,
    240'b101111001111111110111000010100100101010101010101010101010101010101010011010110001010101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111110101110,
    240'b101111001111111110111000010100100101010101010101010101010101010101010101010100110101010010010000111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100111010011111111110101110,
    240'b101111001111111110111000010100100101010101010101010101000101001001010101010101010101010001010000011010111011011011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110001001111001111111111110101110,
    240'b101111001111111110111000010100010101001001001111011010001001111101011101010100110101010101010101010100100101001101110110101100111110010111111101111111111111111111111111111111111111111111111111111100111001001101100010111010111111111110101110,
    240'b101111001111111110110111010110000111001101110011100110101111001101111110010100110101010101010101010101010101010001010001010100100110010010000101101010111100010011010100110111001101101110111111011111010101000001100100111010111111111110101110,
    240'b101111011111111110110100011100101110101111101111111101001111111111000110010101110101010001010101010101010101010101010101010101010101001101010001010100000101010001011011010111110101111101010100010100010101001101100101111010111111111110101110,
    240'b101111011111111110110101011001101110111010110001101000101111001010001001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010001010100010100110101001101010100010101010101001101100101111010111111111110101110,
    240'b101111011111111110111000010011111011110011000010011111001110110001101000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111110111000010011100111101111101010100111011101100001101000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111110111000010100010101011011001111101111000110010101011000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101110111111111110111010010100100101000010001110111010100110100001010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111011011111111010101011,
    240'b101101111111111111011001010110100101000001011101110000001000001101010000010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000100111001111111111110101111010110011010,
    240'b101100011111100111111101101011000110000101011001010111000101110101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110100111001011010110111111111110000010100001,
    240'b110010101101001011111111111111111110010011011010110110101101101011011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111110111111111111111110101011110011011100,
    240'b111100011100011111010111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110000001101000011110011,
    240'b111110001111010111000011101011111011110011000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011011110110010110101111111100011110110,
    240'b111100101111101111010100101101011011011010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011010010110110110111011111001011101111,
    240'b111101001101000011001011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000101110011101101111110011,
    240'b110100101100101011111111111111111111001111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100011101000111010101111101111111111111101001011100111100011,
    240'b101100011111010111111111110000100111010001100111011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001100110011010011000100011100101111111111101100110100110,
    240'b101101101111111111100010011000010100111101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010010010100101001100010010101010100000100110110001010111111011111001110010111,
    240'b101110101111111110111101010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100001001010111101000011001010101000001100110111011111111111010101010,
    240'b101111011111111110111000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110100011100011100111000100110101100101111010111111111110101110,
    240'b101111011111111110111000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000011100010010101111110110010101100101100011111010111111111110101110,
    240'b101111011111111110111000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111100011001110101001110010111001111000011001100000111010111111111110101110,
    240'b101111011111111110111000010100100101010101010101010101010101010001010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101101000001110111001111011110011111100011001100100111010101111111110101110,
    240'b101111011111111110111000010100100101010001010001010100010101010101010100010100010101000001010001010100110101010001010101010101010101010101010101010101010101001001100111111010011111111011110001111101111101101001101100111010011111111110101110,
    240'b101111001111111110111000010100010101010010000001101101011100010011000000101110001010000110000100011001100101010001010001010101000101010101010101010101010101010001011000101100001111011010010100100011010111111001100111111010111111111110101110,
    240'b101111001111111110110111010101001010110011110111111111111111111111111111111111111111111111111100111001111100000110000110010110010101000101010100010101010101010101010001011101101011001001010110010011110100111101100101111010111111111110101110,
    240'b101111001111111110110100100110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111011110011111000001001010100010100100101010101010101010101010101010001010101010101010101001101100101111010111111111110101110,
    240'b101111001111111111000101111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110110011000110101000101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111001111111111100001111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111001101010001010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111001111111111110000111111001111111111111111111111111111111111111111111111111111111111111111111110011101011011010010111010111111111111111111111111111110011001111010010100000101010101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111111101111111111001111111111111111111111111111111111111111111111111111111111111111111101110111111001001111100011011111110111111111111111111111111111100111011101010101000101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111111101010111110111111111111111111111111111111111111111111111111111111111111111111111111111011100001001111010111001101110011111111111111111111111111111111110111010110011001010010010101010101001101100101111010111111111110101110,
    240'b101111011111111111100001111110011111111111111111111111111111111111111111111111111111111111111111111111111110111101101100010011011001111011111111111111111111111111111111111111111100000101010111010101000101001101100101111010111111111110101110,
    240'b101111011111111111010100111101001111111111111111111111111111111111111111111111111111111111111111111111111111111110100110010011100110100011101010111111111111111111111111111111111111110110010101010100000101001101100101111010111111111110101110,
    240'b101111011111111111000111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011000000100111110110011111111111111111111111111111111111111111111100110011001100101000001100101111010111111111110101110,
    240'b101111001111111110111000110010011111111111111111111111111111111111111111111111111111111111101001100100101000101111011000100101000100110001110110111101011111111111111111111111111111111111111111101010010100111101100101111010111111111110101110,
    240'b101111001111111110110011101000101111111111111111111111111111111111111111111111111111111111011110010110010100110111000111110101100101011101010100110001101111111111111111111111111111111111111111111001110110001101100010111010111111111110101110,
    240'b101111001111111110110100011101101111100011111111111111111111111111111111111111111111111111011111010111100101001111000101111111010111111101001011100001101111110011111111111111111111111111111111111111111001010101100000111010111111111110101110,
    240'b101111001111111110110111010101111101011011111111111111111111111111111111111111111111111111011111010111100101001111000100111111111011111001010001010110111101100111111111111111111111111111111111111111111100101001100110111010101111111110101110,
    240'b101111001111111110111000010011011001101011111111111111111111111111111111111111111111111111100011010111100101001111000111111111111111011001110011010011001001100111111111111111111111111111111111111111111110111101111101111010001111111110101110,
    240'b101111001111111110111000010100000110010011100101111111111111111111111111111111111110101010111111010111000101001110101100110110111101110010010001010011110110010111101001111111111111111111111111111111111111110110011110111001101111111110101110,
    240'b101111011111111110111000010100100101000010011100111111111111111111111111111111111010000101010100010101010101010101011001010111000101110001011010010101000101011111011001111111111111111111111111111111111111111111000000111001101111111110101110,
    240'b101111011111111110111000010100100101001101011110110101011111111111111111111111111001100101001001010101010101010101010001010011100100111001001111010011110101001111011000111111111111111111111111111111111111111111011001111010111111111110101110,
    240'b101111011111111110111000010100100101010101010000011111001111010011111111111111111100100110001101010110010101010010000101101000001001111010011110100111101010000011101010111111111111111111111111111111111111111111101100111100011111111110101110,
    240'b101111011111111110111000010100100101010101010101010100011001110111111101111111111111111111100001010111100101001011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101011111111110101110,
    240'b101111011111111110111000010100100101010101010101010101000101010110110010111111111111111111011111010111010101001011000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111101101111111110101110,
    240'b101111001111111110111000010100100101010101010101010101010101001101011000101101111111111111110100110000101011111011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101111111111110101110,
    240'b101111001111111110111000010100100101010101010101010101010101010101010011010110001010101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111110101110,
    240'b101111001111111110111000010100100101010101010101010101010101010101010101010100110101010010010000111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100111010011111111110101110,
    240'b101111001111111110111000010100100101010101010101010101000101001001010101010101010101010001010000011010111011011011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110001001111001111111111110101110,
    240'b101111001111111110111000010100010101001001001111011010001001111101011101010100110101010101010101010100100101001101110110101100111110010111111101111111111111111111111111111111111111111111111111111100111001001101100010111010111111111110101110,
    240'b101111001111111110110111010110000111001101110011100110101111001101111110010100110101010101010101010101010101010001010001010100100110010010000101101010111100010011010100110111001101101110111111011111010101000001100100111010111111111110101110,
    240'b101111011111111110110100011100101110101111101111111101001111111111000110010101110101010001010101010101010101010101010101010101010101001101010001010100000101010001011011010111110101111101010100010100010101001101100101111010111111111110101110,
    240'b101111011111111110110101011001101110111010110001101000101111001010001001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010001010100010100110101001101010100010101010101001101100101111010111111111110101110,
    240'b101111011111111110111000010011111011110011000010011111001110110001101000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111110111000010011100111101111101010100111011101100001101000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101111011111111110111000010100010101011011001111101111000110010101011000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111010111111111110101110,
    240'b101110111111111110111010010100100101000010001110111010100110100001010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101111011011111111010101011,
    240'b101101111111111111011001010110100101000001011101110000001000001101010000010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000100111001111111111110101111010110011010,
    240'b101100011111100111111101101011000110000101011001010111000101110101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110100111001011010110111111111110000010100001,
    240'b110010101101001011111111111111111110010011011010110110101101101011011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111110111111111111111110101011110011011100,
    240'b111100011100011111010111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110000001101000011110011,
    240'b111110001111010111000011101011111011110011000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011011110110010110101111111100011110110,
};
assign data = picture[addr];
endmodule