module Computer();

endmodule