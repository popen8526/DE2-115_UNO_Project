module yellow_three(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110011111011111100001100101101001001110101100101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010111001000010100010111011101111110011111010,
	240'b111111111110100110111011110010111110000011101100111011101110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101110111011001101111111001010110010001111101011111111,
	240'b111110111011101111100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001100011111111110,
	240'b110011001101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110111001110,
	240'b101000101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010011110,
	240'b101010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010101001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000,
	240'b101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
	240'b101000001111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010011110,
	240'b101101111110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010110111,
	240'b111100011011101111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011011111111110101,
	240'b111111101101101010111011111010001111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111100011101111001110101011111110,
	240'b111100101111111111101000101010111010001010101001101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101010101010111010101110101011101010011010000010101000111000111111010011110001,
	240'b111110011111011111100001100101101001001110101100101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010111001000010100010111011101111110011111010,
	240'b111111111110100110111011110010111110000011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111111001010110010001111101011111111,
	240'b111110111011101111100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001100011111111110,
	240'b110011001101010111111111111110101101110011001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111011001101110011101101111111111100111111111100110111001110,
	240'b101000101111100011111110110010111010100010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001101010111010111010101011001010100011010011111111111110111010011110,
	240'b101010001111111111110001101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100101110101011111011111001011010110110110011111110001111110110101001,
	240'b101011101111111111101011101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110010001111011011001010111001101011100110101110111100101111111110110000,
	240'b101011101111111111101011101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110000101111100011011001101101011010100110110000111100101111111110110000,
	240'b101011101111111111101011101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110011101111110111110000101101111010011110110000111100101111111110110000,
	240'b101011101111111111101011101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101110111100001101011110101101101010111010101110110000111100101111111110110000,
	240'b101011101111111111101011101011001010100110101001101010001010011110101000101010001010100010101001101010101010101010101010101010101010101010101010101010101010100110110001111101011100011010100010110010011101110010110010111100101111111110110000,
	240'b101011101111111111101011101011001010011110101110110000011100110011001011110001111011110010110010101010101010100010101001101010101010101010101010101010101010101010101010111000101111001011010110111101111101101010101111111100101111111110110001,
	240'b101011101111111111101011101010111011101011101001111111101111111111111111111111111111110011110011111000111100110010110100101010011010100010101010101010101010101010101001101101011110010011110011110111101011000010101111111100101111111110110001,
	240'b101011101111111111101001101110011111000111111111111111111111111111111111111111111111111111111111111111111111111111110101110110001011010110101000101010011010101010101010101010011010101110110000101010101010100010110000111100101111111110110001,
	240'b101011101111111111101010110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011001101101010111010100110101010101010101010101010101001101010101010100110110000111100101111111110110001,
	240'b101011101111111111110001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011011001010101000101010101010101010101010101010101010100110110000111100101111111110110001,
	240'b101011101111111111111000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110011111111111111111111111111110101110110110101010001010101010101010101010101010100110110000111100101111111110110001,
	240'b101011101111111111111001111111001111111111111111111111111111111111111111111111111111111111111111111101101100110010111000101110001101000011111001111111111111111111101110101101101010100010101010101010101010100110110000111100101111111110110000,
	240'b101011101111111111110111111110111111111111111111111111111111111111111111111111111111111111111001110000001010011010100111101001111010011111000111111111001111111111111111111010101011000010101001101010101010100110110000111100101111111110110000,
	240'b101011101111111111110100111110011111111111111111111111111111111111111111111111111111111111011101101010001010101010111010101101111010100010101001111001011111111111111111111111111101110110101010101010101010100110110000111100101111111110110000,
	240'b101011101111111111110000111101011111111111111111111111111111111111111111111111111111111111001010101001011011100111111000111100101011100010101101110101101111111111111111111111111111110111001000101010001010100110110000111100101111111110110000,
	240'b101011101111111111101100111010101111111111111111111111111111111111111111111111111111111111001000101001011011110011111100111111111111010011101111111101101111111111111111111111111111111111110010101100101010100010110000111100101111111110110000,
	240'b101011101111111111101000110110101111111111111111111111111111111111111111111111111111111111011001101010001010101111000100110100001110110111111111111111111111111111111111111111111111111111111111110101001010011110110000111100101111111110110001,
	240'b101011101111111111101000110010001111111011111111111111111111111111111111111111111111111111101010101011011010100110101000101001101101101111111111111111111111111111111111111111111111111111111111111101001011001010101111111100101111111110110001,
	240'b101011101111111111101001101101011111010011111111111111111111111111111111111111111111101011000000101010011010100010101010101011001101110111111111111111111111111111111111111111111111111111111111111111111100110010101110111100101111111110110001,
	240'b101011101111111111101010101010111101111011111111111111111111111111111111111111111101110010101000101010011100010111100111111011001111011111111111111111111111111111111111111111111111111111111111111111111110011110110001111100101111111110110001,
	240'b101011101111111111101011101010101100000011111101111111111111111111111111111111111100001010100101101110101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110111110111100001111111110110001,
	240'b101011101111111111101011101011001010101111100111111111111111111111111111111110111011100110100101110100001111111111111111111111111111111111110101111011101111001111111111111111111111111111111111111111111111111111010000111011111111111110110000,
	240'b101011101111111111101011101011001010011111000001111111001111111111111111111111001011101010100101110011001111111111111111111111111111111111000110101010011100010011111111111111111111111111111111111111111111111111100001111100001111111110110000,
	240'b101011101111111111101011101011001010100110101010110111101111111111111111111111111100011110100110101101001111000111111111111111111110101010101111101001011101000011111111111111111111111111111111111111111111111111101110111100111111111110110000,
	240'b101011101111111111101011101011001010100110101000101100111111001011111111111111111110010110101010101010001011100011011000110101011011010010101000101011011110110011111111111111111111111111111111111111111111111111110111111101101111111110110000,
	240'b101011101111111111101011101011001010100110101010101010001100001011111010111111111111110111001100101010001010011110100111101001111010011110101001110101001111111111111111111111111111111111111111111111111111111111111100111110001111111110110000,
	240'b101011101111111111101011101011001010100110101010101010101010100011001101111111011111111111111011110100011011001010101001101010101011010011010111111111011111111111111111111111111111111111111111111111111111111111111100111110011111111110110000,
	240'b101011101111111111101011101011001010100110101010101010101010101010101001110011111111110011111111111111111111001011100110111001111111010011111111111111111111111111111111111111111111111111111111111111111111111111111100111110101111111110110001,
	240'b101011101111111111101011101011001010100110101010101010101010101010101001101010011100100111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101111111111110110001,
	240'b101011101111111111101011101011001010100110101010101010101010101010101010101010101010100010111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101111100101111111110110001,
	240'b101011101111111111101011101011001010100110101000101010001010100010101010101010101010101010101000101011101100110011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000001111100001111111110110001,
	240'b101011101111111111101011101011001010101111001010110111011100011010101010101010101010101010101010101010011010100010110010110010101110011111111001111111111111111111111111111111111111111111111111111101101100010110101110111100101111111110110001,
	240'b101011101111111111101011101010111101001011111011111011101111101011001011101010001010101010101010101010101010101010101001101010001010110010111000110010001101011111100000111001011110010111010111101110011010011110110000111100101111111110110000,
	240'b101011101111111111101010101100011110101111010001101010101101101111101011101011001010100110101010101010101010101010101010101010101010100110101000101010001010100010101001101010111010101010101000101010001010100110110000111100101111111110110000,
	240'b101011101111111111101011101011101011011010101101101001011101001111101110101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111100101111111110110000,
	240'b101011101111111111101011101011001010011110111000110111101111011111010100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111100101111111110110000,
	240'b101011101111111111101011101011001010011110111011111100011111100110111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111100101111111110110000,
	240'b101011101111111111101011101010111011100111010000101111111111100111000001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111100101111111110110000,
	240'b101010111111111111101101101010111011101011111000111101011111001010110101101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110001111101011111111110101110,
	240'b101000001111110111111010101111001010010110111110110101001011101110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011011000100111111101111010010011110,
	240'b101101111110001011111111111011101100001110111000101110001011100110111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100011111110011111111111101101010110111,
	240'b111100011011101111110110111111111111111011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111100011011111111110101,
	240'b111111101101101010111011111010001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100011101111001110101011111110,
	240'b111100101111111111101000101010111010001010101001101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101010101010111010101110101011101010011010000010101000111000111111010011110001,
	240'b111110011111011111100001100101101001001110101100101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010111001000010100010111011101111110011111010,
	240'b111111111110100110111011110010111110000111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111111001010110010001111101011111111,
	240'b111110111011101111100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001100011111111110,
	240'b110011001101010111111111111100011001011001101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110110101101001011011101010000011110111111111111100110111001110,
	240'b101000101111100111111011011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110000000001100000000001111011111111101110111110011110,
	240'b101010001111111111010100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011100000011110100101100000000110000011010111010001111111010101001,
	240'b101011101111111111000001000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110111110010001100000101100110010110000001101110110001111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111110110010001100001000010000001100010011110110001111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011001111100111010010001001010000000000010011110110001111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110110100111000011100001111000000100000010100010100110110001111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101111000100101010100000000010111101001011100010111110101111111111110110000,
	240'b101011101111111111000010000010000000000000001100010001100110011001100100010101100011010100011001000000000000000000000000000000000000000000000000000000000000000000000100101010001101100110000100111010001000111000001110110110001111111110110001,
	240'b101011101111111111000010000000100011001010111110111110111111111111111111111111101111011111011011101011000110011000011111000000000000000000000000000000000000000000000000001000011010110111011010100111010001001000010000110110001111111110110001,
	240'b101011101111111110111101001011011101011111111111111111111111111111111111111111111111111111111111111111111111111111100000100010110010001100000000000000000000000000000000000000000000001100010011000000000000000000010011110110001111111110110001,
	240'b101011101111111110111111101000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101101001000001100000000000000000000000000000000000000000000000000000000000010011110110001111111110110001,
	240'b101011101111111111010110111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001000001100100000000000000000000000000000000000000000000000000010011110110001111111110110001,
	240'b101011101111111111101000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111011011111111111111111111111111100001100100110000000000000000000000000000000000000000000010011110110001111111110110001,
	240'b101011101111111111101011111101011111111111111111111111111111111111111111111111111111111111111111111000110110011000101010001011000111010011101100111111111111111111001100001001010000000000000000000000000000000000010011110110001111111110110000,
	240'b101011101111111111100110111100101111111111111111111111111111111111111111111111111111111111101110010000110000000000000000000000000000000001011000111101101111111111111111110000010001010100000000000000000000000000010011110110001111111110110000,
	240'b101011101111111111011101111011101111111111111111111111111111111111111111111111111111111110011001000000000000000000101111001010000000000000000000101100011111111111111111111111111001100100000100000000000000000000010011110110001111111110110000,
	240'b101011101111111111010000111000011111111111111111111111111111111111111111111111111111111101011111000000000010101111101010110110000010101000001110100001011111111111111111111111111111101101011010000000000000000000010011110110001111111110110000,
	240'b101011101111111111000101110000011111111111111111111111111111111111111111111111111111111101011010000000000011010111111000111111111101110111001111111001011111111111111111111111111111111111010111000110010000000000010011110110001111111110110000,
	240'b101011101111111110111010100100011111111111111111111111111111111111111111111111111111111110001111000000010000010001001110011100011100100111111111111111111111111111111111111111111111111111111111011111100000000000010011110110001111111110110001,
	240'b101011101111111110111010010110011111110111111111111111111111111111111111111111111111111111000010000010100000000000000000000000001001001111111111111111111111111111111111111111111111111111111111110111100001011100001111110110001111111110110001,
	240'b101011101111111110111110001000011101111011111111111111111111111111111111111111111110111101000010000000000000000000000001000010001001101111111111111111111111111111111111111111111111111111111111111111110110010100001011110110001111111110110001,
	240'b101011101111111111000001000001001001110111111111111111111111111111111111111111111001011100000000000000000101000010110110110001101110100011111111111111111111111111111111111111111111111111111111111111111011011100010111110101111111111110110001,
	240'b101011101111111111000010000000010100000011111000111111111111111111111111111111010100100100000000001100011110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101100111101110100111111111110110001,
	240'b101011101111111111000010000001100000011010111000111111111111111111111111111100100010110100000000011100011111111111111111111111111111111111100010110011001101101011111111111111111111111111111111111111111111111101110010110100001111111110110000,
	240'b101011101111111111000010000010000000000001000101111101111111111111111111111101010011000100000000011010001111111111111111111111111111111101010101000010010100111111111111111111111111111111111111111111111111111110100110110100101111111110110000,
	240'b101011101111111111000010000010000000000000000011100110111111111111111111111111110101100000000000000111111101010011111111111111111100001000010001000000000111001011111111111111111111111111111111111111111111111111001100110111001111111110110000,
	240'b101011101111111111000010000010000000000000000000000111011101011111111111111111111011000000000011000000000010101010001000100000010001111100000000000011001100011111111111111111111111111111111111111111111111111111101000111001011111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000100011111101111111111111111101001100111000000000000000000000000000000000000000000000000011111111111111011111111111111111111111111111111111111111111111111110101111010111111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000000000001101000111110001111111111110011011101100001100100000000000000000001111010001000111110011111111111111111111111111111111111111111111111111111111111110110111011101111111110110000,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000011011111111011111111111111111111101100110110101101101111101111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011101111111110110001,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000101110011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111001111111111110110001,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000000000000110110101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000110101101111111110110001,
	240'b101011101111111111000010000010000000000000000000000000000000000000000000000000000000000000000000000011000110100011010011111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101000110110100111111111110110001,
	240'b101011101111111111000010000001100000010101100000100110000101010100000011000000000000000000000000000000000000000000011001011000011011100111101100111111111111111111111111111111111111111111111111111001000101000100001110110110001111111110110001,
	240'b101011101111111111000001000000110111100111110010110011001111001001100010000000000000000000000000000000000000000000000000000000000000011000101011010110111000010110100011101011111011000010000110001011000000000000010010110110001111111110110000,
	240'b101011101111111110111111000101011100010001110111000010101001001111000101000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000010011110110001111111110110000,
	240'b101011101111111111000001000011010010010000001000000000000111110011001011000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110001111111110110000,
	240'b101011101111111111000010000010000000000000101010100110111110100001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110001111111110110000,
	240'b101011101111111111000010000010000000000000110100110101011110111000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110001111111110110000,
	240'b101011101111111111000001000000110010111001110010001111111110101101000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110001111111110110000,
	240'b101010111111111111001010000001000011000011101010111000101101100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101111000001111111110101110,
	240'b101000001111110111110001001101110000000000111101011111100011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001110111110101111010110011110,
	240'b101101111110001011111111110011000100111000101010001010110010110000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000101100011011010111111111101101010110111,
	240'b111100011011101111110110111111111111101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101111110111111111111100011011111111110101,
	240'b111111101101101010111011111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100011101111001110101011111110,
	240'b111100101111111111101000101010111010001010101001101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101010101010111010101110101011101010011010000010101000111000111111010011110001,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule