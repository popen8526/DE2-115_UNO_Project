module yellow_skip(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110101111110011101011101000101000111110101010101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010011000110110101100111100111111110011111010,
	240'b111111111111101111000010110001101101111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010111101110111000111110011101111110111111111,
	240'b111111111100110011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101000111111110,
	240'b110011011100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011111001100,
	240'b100111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010010011010,
	240'b101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110101111,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011000000,
	240'b101100101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110110101,
	240'b100111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010011010,
	240'b101111001101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101110111100,
	240'b111110111100010011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011100100011111001,
	240'b111111011111000110111100110110011111011011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111010111010101110000001111010111111101,
	240'b111100001111001111110100101100001001110010101001101010111010101010101010101010101010101010101010101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001101010101100111011001111001011110000,
	240'b111110101111110011101011101000101000111110101010101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010011000110110101100111100111111110011111010,
	240'b111111111111101111000010110001101101111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010111101110111000111110011101111110111111111,
	240'b111111111100110011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101000111111110,
	240'b110011011100101011111111111111011110000011001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001110110011011100110011001110110011111110001111111110111111101100011111001100,
	240'b100111111110011111111111110101101010100110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011010101001101110001011101110101101101001011010101011011100111111111110010110011010,
	240'b101011111111100011111011101101111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011010011100100111110001111101011101111110000011010010110111100111111011111000010101111,
	240'b101101101111110011110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011001110011011111111110100001011110111100011111101101011010110110101111110101110111111000000,
	240'b101101101111110011110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110000001111100011110011111001101010110010101011111011101101010110110100111110101110111111000000,
	240'b101101101111110011110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110100001110101010111011111101001110001010101001110101101110010110110111111110101110111111000000,
	240'b101101101111110011110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110011011110111110101010101111011111100011011000110111011110001010110110111110101110111111000000,
	240'b101101101111110011110110101100111010100110101001101010001010100010101000101010001010100010101001101010101010101010101010101010101010101010101000101110101111100111001000101001001100001011111001111111101100110010110100111110101110111111000000,
	240'b101101111111110011110110101100111010011110101100110000001100110111001101110010011011111110110100101010111010100010101000101010101010101010101010101010011101011111111010110111001101011011111010111010101010111010110110111110101111000011000000,
	240'b101101111111110011110110101100011011010111100101111111011111111111111111111111111111111011110101111001101100111110110110101010011010100010101010101010011010110011010000111011101111000011011011101100111010011110110111111110101111000011000000,
	240'b101101111111110011110100101110011110101011111111111111111111111111111111111111111111111111111111111111111111111111110110110110111011011110101000101010011010100110101000101011011010111010101001101010011010100010110111111110101111000011000000,
	240'b101101111111110011110011110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011001110101011001010100110101010101010011010100110101010101010101010100010110111111110101111000011000000,
	240'b101101111111101111110111111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101011001010101000101010101010101010101010101010101010100010110111111110101111000011000000,
	240'b101101101111101111111010111111001111111111111111111111111111111111111111111111111111111111111111111111111111110011110110111101101111110011111111111111111110101110110110101010001010101010101010101010101010100010110111111110101110111111000000,
	240'b101101101111101111111010111111001111111111111111111111111111111111111111111111111111111111110100110101001011110010110101101101011011110111010110111101101111111111101101101101011010100010101010101010101010100010110111111110101110111111000000,
	240'b101101101111101111111010111110111111111111111111111111111111111111111111111111111110010110110110101001111010011010100110101001101010011110101000101110001110100111111111111010001010111110101001101010101010100010110111111110101110111111000000,
	240'b101101101111101111111000111110001111111111111111111111111111111111111111111001111010111110101000101010111011011011000011110000101011010010101000101001111011001011101011111111111101101010101001101010101010100010110111111110101110111111000000,
	240'b101101101111101111110110111011111111111111111111111111111111111111110110101110001010100010101000101110101111010011111111111111101111010111010001101010111010011110111011111110011111110111000100101010001010100010110111111110101110111111000000,
	240'b101101101111110011110100111000111111111111111111111111111111111111010111101001111010100110101000101010111101011111111111111111111111111111111111110101001010100110101000110111011111111111101110101011111010011110110111111110101110111111000000,
	240'b101101111111110011110011110100111111111111111111111111111111110010111101101001101011100110110110101001111010101111011110111111111111111111111111111110101011101110100110110000011111111011111111110011101010011010110111111110101111000011000000,
	240'b101101111111110011110100110000101111100111111111111111111111001010110000101001111101110111101100101100011010011110101110111001011111111111111111111111111101011010100110101100111111011011111111111011111010110110110110111110101111000011000000,
	240'b101101111111110011110101101101011110100111111111111111111110110010101010101010101110101111111111111000111010110110100111101100101110101111111111111111111110010010101001101011101110111111111111111111101100010010110100111110101111000011000000,
	240'b101101111111110011110101101100001101000011111111111111111110101110101010101010101110110011111111111111111101110010101011101001111011011111110001111111111110010110101001101011101110111011111111111111111101111110110110111110101111000011000000,
	240'b101101111111110011110110101100011011010011110111111111111111000110101110101010001110000111111111111111111111111111010101101010011010011110111100111101111101110010100111101100011111010011111111111111111111001111000000111110011111000011000000,
	240'b101101101111110011110110101100111010011111011010111111111111101010111001101001101100011111111111111111111111111111111101110011011010100010100111110000111011111010100110101111011111110011111111111111111111110111001110111110001110111111000000,
	240'b101101101111110011110110101100111010011110110111111101111111111111010001101001111010110011100100111111111111111111111111111110111100011110101001101010011010100110101000110101101111111111111111111111111111111111011110111110001110111111000000,
	240'b101101101111110011110110101100111010100110101000110100011111111111110001101100101010011110110011111001001111110111111111111111111111010010110110101010001010100010110101111101011111111111111111111111111111111111101100111110001110111111000000,
	240'b101101101111110011110110101100111010100110101001101011011110100011111111110111001010101010100111101011011100001011010011110100101100000110101101101010001010110011100001111111111111111111111111111111111111111111110100111110101110111111000000,
	240'b101101101111110011110110101100111010100110101010101010001011100011110100111111111101011110101101101001111010011110100111101001111010011110100111101011111101110011111111111111111111111111111111111111111111111111110111111111001110111111000000,
	240'b101101101111110011110110101100111010100110101010101010101010100011000010111110011111111111100111110000111011000110101010101010101011001011000110111010111111111111111111111111111111111111111111111111111111111111111000111111011110111111000000,
	240'b101101111111110011110110101100111010100110101010101010101010101010101000110001011111100011111111111111101111001011101010111010101111001111111111111111111111111111111111111111111111111111111111111111111111111111111001111111011110111111000000,
	240'b101101111111110011110110101100111010100110101010101010101010101010101010101010001100000011110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111110101110111111000000,
	240'b101101111111110011110110101100111010100110101010101010101010101010101010101010101010100010110101111000001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111110001110111111000000,
	240'b101101111111110011110110101100111010100110101001101010001010100110101001101010001010101010101000101010111100010111101011111111101111111111111111111111111111111111111111111111111111111111111111111111111110111010111111111110011111000011000000,
	240'b101101111111110011110110101100111010100010101110110011011110001111011101101111101010100110101010101010011010100010101110110001001110001011110101111111101111111111111111111111111111111111111111111011101011101010110101111110101111000011000000,
	240'b101101101111110011110110101100101010110011100010111110111110011011101101111110011100011010101000101010101010101010101001101010001010101010110100110000111101000011011010110111111101111011001110101100101010011110110111111110101110111111000000,
	240'b101101101111110011110101101100001100101011111111111101011011100010101011110110101111001110110010101010011010101010101010101010101010101010101001101010001010011110101000101010011010100110100111101010011010100010110111111110101110111111000000,
	240'b101101101111110011110101101100101110010111100001111010101110110110110000101100001111010111000100101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110111111110101110111111000000,
	240'b101101101111110011110101101101001110101111001101101100111111001011100110101100011111000011001011101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110111111110101110111111000000,
	240'b101101101111110011110101101100011110000111100001101001011011101011110101111010001111010111000000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110111111110101110111111000000,
	240'b101101111111110011110101101100001100001011111010110011101010111111001111111111111110101010101101101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110111111110101110111111000000,
	240'b101100101111101011111001101101001010100011010011111110101111010111111000111011101011101010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111111001111000010110101,
	240'b100111111110101111111111110011001010011010100111101110101100110011000111101011111010011010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011111010010111111111110100110011010,
	240'b101111001101000111111111111110001101000011000000101111111011111010111110101111111100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001101001111111010111111111100101110111100,
	240'b111110111100010011100110111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111111111000011100100011111001,
	240'b111111011111000110111100110110011111011111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111011011010101110000001111010111111101,
	240'b111100001111001111110100101100001001110010101001101010111010101010101010101010101010101010101010101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001101010101100111011001111001011110000,
	240'b111110101111110011101011101000101000111110101010101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010011000110110101100111100111111110011111010,
	240'b111111111111101111000010110001101101111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010111101110111000111110011101111110111111111,
	240'b111111111100110011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101000111111110,
	240'b110011011100101011111111111110001010001001101111011011010110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101100011010000110011101101010011100001010101011111011111111101100011111001100,
	240'b100111111110100011111111100001010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110011001100001010000000000000010010010101111111111110010110011010,
	240'b101011111111101011110000001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110101110111010101110111111010000010001010000000000110101111101101111000110101111,
	240'b101101101111111011100010000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011011010011111111011100010011111110101011111000100010001100100010111011011111000111000000,
	240'b101101101111111011100010000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111110101011011011101101010000101100001001110010101000001000100000111011011111001011000000,
	240'b101101101111111011100010000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111100000000110010110111011010100000000100100001001011000000100111111011001111001011000000,
	240'b101101101111111011100010000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010101100111000000001001110101110101010001010100110001010100000100110111011001111001011000000,
	240'b101101101111111011100010000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111110101101011011000000000100100111101100111110110110010100011111111011011111001011000000,
	240'b101101111111111011100010000110110000000000001000010000110110101101101010010111100011110100011111000000100000000000000000000000000000000000000000000000011000011111110000100101111000010111110000110000100000111100100100111011011111001011000000,
	240'b101101111111111011100010000101100010001010110010111110101111111111111111111111111111101111100010101101010111000000100101000000000000000000000000000000000000011101110000110010111101001010010011000110110000000000100111111011011111001011000000,
	240'b101101111111111011011111001011101100000011111111111111111111111111111111111111111111111111111111111111111111111111100101100100110010100000000000000000000000000000000000000010010000111000000000000000000000000000100111111011011111001011000000,
	240'b101101111111111011011011100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001101101101000001110000000000000000000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101111111110111100110110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010000001101000000000000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101101111110011101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111011011100011111000111111011111111111111111111100001100100101000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101101111110011110000111101011111111111111111111111111111111111111111111111111111111111011101011111100011100000100010001000100011101010000100111000111111111111001010001000100000000000000000000000000000000000100111111011011111001011000000,
	240'b101101101111110011101110111101001111111111111111111111111111111111111111111111111011000000100100000000000000000000000000000000000000000000000000001010111011110011111111101110110001000100000000000000000000000000100111111011011111001011000000,
	240'b101101101111110011101010111010101111111111111111111111111111111111111111101101110001000100000000000000110010010101001101010010000001111100000000000000000001100111000100111111111001000000000001000000000000000000100111111011011111001011000000,
	240'b101101101111110111100100110011111111111111111111111111111111111111100101001010010000000000000000001100001101111111111110111111011110000001110101000001110000000000110100111011101111100001001110000000000000000000100111111011011111001011000000,
	240'b101101101111111011011100101010111111111111111111111111111111111110000111000000000000000000000000000001111000011111111111111111111111111111111111100000000000000100000000100110001111111111001100000100010000000000100111111011011111001011000000,
	240'b101101111111111011011010011110101111111011111111111111111111011000111000000000000010111000100100000000000000011110011010111111111111111111111111111100100011010000000000010001101111101111111111011011010000000000100111111011011111001011000000,
	240'b101101111111111011011101010010001110110111111111111111111101100100010010000000001001101011000101000101100000000000001111101100001111111111111111111111111000010100000000000110101110011011111111110100000000110000100100111011011111001011000000,
	240'b101101111111111011100000001000011011110111111111111111111100011000000010000000001100001011111111101010100000110000000000000110011100001111111111111111111010111100000000000011001101000011111111111111010100111100011111111011011111001011000000,
	240'b101101111111111011100010000100110111000111111111111111111100010000000001000000011100011011111111111111111001010100000110000000000010011111010100111111111011001000000000000011001100111011111111111111111001111100100100111011001111001011000000,
	240'b101101111111111011100010000101100001111111101000111111111101010000001100000000001010001111111111111111111111111001111111000000010000000000111000111010001001010100000000000101011110000011111111111111111101110001000001111010011111001011000000,
	240'b101101101111111011100010000110100000000010010010111111111111000000101101000000000101011011111110111111111111111111111001011010010000000000000000010010110011111000000000001110011111011111111111111111111111100001101101111001101111001011000000,
	240'b101101101111111011100010000110110000000000100110111001111111111101110100000000000000100110101110111111111111111111111111111100110101100000000000000000000000000000000000100001001111111111111111111111111111111110011110111001101111000111000000,
	240'b101101101111111011100010000110110000000000000000011101101111111111010110000101110000000000011100101011111111101011111111111111111101111000100100000000000000000000100001111000001111111111111111111111111111111111000111111001111111000111000000,
	240'b101101101111111011100010000110110000000000000000000011001011101111111111100101010000001100000000000010000100100101111100011110000100010000001010000000000000100010100110111111111111111111111111111111111111111111011101111011001111000111000000,
	240'b101101101111111011100010000110110000000000000000000000000010101111011111111111111000011100001010000000000000000000000000000000000000000000000000000100011001011011111111111111111111111111111111111111111111111111100111111100101111000011000000,
	240'b101101101111111011100010000110110000000000000000000000000000000001001001111011001111111110111000010011000001010100000001000000010001100101010100110000111111111111111111111111111111111111111111111111111111111111101100111101011111000011000000,
	240'b101101111111111011100010000110110000000000000000000000000000000000000000010100011110101111111111111110111101011111000000110000001101101111111110111111111111111111111111111111111111111111111111111111111111111111101100111101011111000011000000,
	240'b101101111111111011100010000110110000000000000000000000000000000000000000000000000100001011011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111011011111000011000000,
	240'b101101111111111011100010000110110000000000000000000000000000000000000000000000000000000000100100101000111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000111001101111000111000000,
	240'b101101111111111011100010000110110000000000000000000000000000000000000000000000000000000000000000000001000101001111000011111111011111111111111111111111111111111111111111111111111111111111111111111111111100110001000000111010011111001011000000,
	240'b101101111111111011100010000110110000000000001100011010101010110010011001001111000000000000000000000000000000000000001110010100001010011111100010111110111111111111111111111111111111111111111111110011010011000000100010111011011111001011000000,
	240'b101101101111111011100010000110000000100110101000111100101011010011001001111011100101011000000000000000000000000000000000000000000000000100011110010010100111001110010000100111101001101101101100000110000000000000100111111011011111001011000000,
	240'b101101101111111011100010000101000101111111111111111000100010101000001000100100001101101100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101101111111011100001000110011011000010100101101111101100100000010100000100111110000001001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101101111111011100000000111111100010001101010000111011101100110110100000101001101000101100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101101111111011100001000101101010011010100101000000000011000011011111101110001110001001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111011011111001011000000,
	240'b101101111111111011100010000101000100100011110001011011000001011001110000111111111100000000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110111011011111001011000000,
	240'b101100101111110011101011000111100000000001111011111100001110000111101010110011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111100111111000110110101,
	240'b100111111110110011111110011001110000000000000000001100000110100001010110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111111111111110100110011010,
	240'b101111001101000111111111111010100111001101000010001111010011110000111100010000000100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010001000111101111110000111111111100101110111100,
	240'b111110111100010011100110111111111111111111111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110011111111111111111111000011100100011111001,
	240'b111111011111000110111100110110011111011111111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111011011010101110000001111010111111101,
	240'b111100001111001111110100101100001001110010101001101010111010101010101010101010101010101010101010101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001101010101100111011001111001011110000,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule