module red_eight(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111011111111001111110000110001111011000110110010101100111011001010110010101100101011001010110011101100111011001110110011101100111011001110110010101100101011001010110010101100111011001110110011101100111011000110111011111000011111001011101111,
	240'b111100011110100011000000110110001111011111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111100001101110011101101011110010,
	240'b111010101011110011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011101111100100,
	240'b101100101101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001110110011,
	240'b100100101110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011011,
	240'b101010011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101,
	240'b101011011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100,
	240'b100101011111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100,
	240'b101010001101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101011,
	240'b111001011011101111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111011011101,
	240'b111100101110000010111101111010001111111111111110111111011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011110001101111111101000011110010,
	240'b111110011111101111100101101001011001011010101110101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001001110010011101110111101111110011111001,
	240'b111011111111001111110001110001111011001010110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011000110111100111000011111001011101111,
	240'b111100011110100011000000110110001111011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101011100001101110011101101011110010,
	240'b111010101011110011101000111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111111111111111111101001011101111100100,
	240'b101100101101000111111111111100011010010001111110011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111101101111000011110101001010111100011111111111110001110110011,
	240'b100100101110111011111110100110110100111001010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110110011110010100011100110100101101111100111101011111111010011011,
	240'b101010011111100111110011011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011000011101011111110100111010100111001101010101110101111111111110110000,
	240'b101101011111101111101101011000110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011111001111000010001100111001111001101001010001110100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011011001110110111011101111101101000010101010001110100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100101001111010111010100111100011011001001010100110100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100111011101001010000100101111110100001100110110011101111111110111100,
	240'b101101011111101111101101011001000101001101010011010100000101000101010010010100000100111101010001010100110101010001010101010101010101010101010101010101010101010001010111110101101011001101001100100100011110101001101000110011101111111110111100,
	240'b101101011111101111101101011001000100111101100010100101001010111110110000101010001001011101111110011000110101010001010000010101000101010101010101010101010101010101010001100111111111011011000111111011111011110101010110110100001111111110111100,
	240'b101101011111101111101101011000000111011011011010111111111111111111111111111111111111111111111001111001101011111110001001010110110101000001010100010101010101010101010100010110101010001011010010101100100110001101010100110100001111111110111100,
	240'b101101011111101111101010011101111110000011111111111111111111111111111111111111111111111111111111111111111111111111111100110101001000101101010110010100100101010101010101010101000101001001010111010100110101001001010110110100001111111110111100,
	240'b101101011111101111101001101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111000010011010110101000101010101010101010101010101010100010101010101010001010110110100001111111110111100,
	240'b101101011111100111110011111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011000001101010001010101000101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111100111111010111111001111111111111111111111111111111111111111111111111111111111111111111111111111111011101010111001111111101011111111111111111111001010001111010100010101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111100111111011111111011111111111111111111111111111111111111111111111111111111111111111111011101001010101100010010111111000001111011101111111111111111111110100100010110101000001010101010101010101010001010110110100001111111110111100,
	240'b101101011111100111111001111110001111111111111111111111111111111111111111111111111111111111111000100010110100111001001111010011100100111001110001111010101111111111111111111011110111100101010001010101010101010001010110110100001111111110111100,
	240'b101101011111100111110101111011011111111111111111111111111111111111111111111111111111111111001111010101010101001101111001100001000101011101001111101011011111111111111111111111111101101101100011010100110101010001010110110100001111111110111100,
	240'b101101011111101011101111110110111111111111111111111111111111111111111111111111111111111110101100010011100110010111100111111111000111110001001100100010111111111011111111111111111111111110110100010100110101010001010110110100001111111110111100,
	240'b101101011111101111101001110001001111111111111111111111111111111111111111111111111111111110101100010011100110010111100110111110100111101101001100100010111111111011111111111111111111111111110111011111010101000001010110110100001111111110111100,
	240'b101101011111101111101000101000101111111111111111111111111111111111111111111111111111111111010011010110100101001101110110100000010101011101010001101100011111111111111111111111111111111111111111110010010101011001010101110100001111111110111100,
	240'b101101011111101111101010100000011111001011111111111111111111111111111111111111111111111111100111011001110101001001010000010011110101001101011000110010111111111111111111111111111111111111111111111110010111110001010010110100001111111110111100,
	240'b101101011111101111101100011001111101000111111111111111111111111111111111111111111111101010001111010100100101001001011010010111010101001101010001011101011110110111111111111111111111111111111111111111111011100101010011110100001111111110111100,
	240'b101101011111101111101101010111111001111011111111111111111111111111111111111111111100110101010110010100011000001011010011110111001001101001010101010011111010110011111111111111111111111111111111111111111110100001100110110011101111111110111100,
	240'b101101011111101111101101011000010110100011101110111111111111111111111111111111111001110101001101011010001110100011111111111111111111101010000000010011000111110011111010111111111111111111111111111111111111110110001011110010111111111110111100,
	240'b101101011111101111101101011001000101000010110011111111111111111111111111111111111000100101001011100010011111111111111111111111111111111110101010010011010110110111110000111111111111111111111111111111111111111110110010110010111111111110111100,
	240'b101101011111101111101101011001000100111101101100111011011111111111111111111111111000111001001011100000011111110111111111111111111111111110100001010011000111000111110011111111111111111111111111111111111111111111010011110100111111111110111100,
	240'b101101011111101111101101011001000101001101010001101000001111111111111111111111111010110101001110010111001100110011111111111111111110010001101100010011011000100111111110111111111111111111111111111111111111111111101001110110111111111110111100,
	240'b101101011111101111101101011001000101001101010011010110101100111011111111111111111110001001100001010100000110010110100001101010010111000101010001010101001100010111111111111111111111111111111111111111111111111111110010111001111111111110111100,
	240'b101101011111101111101101011001000101001101010101010100010110111011100101111111111111111110110100010101010100111101010000010100000100111101010000100101011111101011111111111111111111111111111111111111111111111111110111111100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101000010000000111011101111111111111101101110010110111001010111010101110110010110100011111101101111111111111111111111111111111111111111111111111111111111111001111101011111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010000100001011110111011111111111111111110111111010010110011101110100011111111111111111111111111111111111111111111111111111111111111111111111111111010111101101111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010100010111110111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111010101111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101000001101100110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000110101011111111110111100,
	240'b101101011111101111101101011001000101001001010001010100100101000101010100010101010101010101010010010101111000111011011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001110110011001111111110111100,
	240'b101101011111101111101101011001000101001010001000101101101001100101011011010101000101010101010101010101000101000001011111100100001100101111110000111111101111111111111111111111111111111111111111111101101010001001010101110100001111111110111100,
	240'b101101011111101111101101011000001000101011110101111000101111011110101101010100110101010101010101010101010101010101010011010100000101011101101101100011111010101111000000110010111100111010111000011111100101001001010101110100001111111110111100,
	240'b101101011111101111101101011000111100111111000000010101101001110011101100011000110101001101010101010101010101010101010101010101010101010001010010010100000101000001010100010101110101100001010011010100010101010001010110110100001111111110111100,
	240'b101101011111101111101100011001001101011010110000010010001000100011110000011001100101001101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001010110110100001111111110111100,
	240'b101101011111101111101101011000001001111011110000101110011110010011000011010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111101111101101011000010110011111101110111100101111101110000111010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111101111101101011000000111100011101110100010101110000110011110010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100001111111110111101,
	240'b101011011111101011110001011001000110001111100010111001101111000101111111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110101001111111110110100,
	240'b100101011111000111111101100011010100101101111000101101101000110001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100111001110000111100001111111110011100,
	240'b101010001101100011111111111001101000100101100111011001100110011101101010011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010100111110011010010111111111110101010101011,
	240'b111001011011101111110001111111111111101111110001111100001111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100001111100011111111111110111011111011011101,
	240'b111100101110000010111101111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001101111111101000011110010,
	240'b111110011111101111100101101001011001011010101110101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001001110010011101110111101111110011111001,
	240'b111011111111001111110000110001111011000110110010101100111011001010110010101100101011001010110011101100111011001110110011101100111011001110110010101100101011001010110010101100111011001110110011101100111011000110111011111000011111001011101111,
	240'b111100011110100011000000110110001111011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101011100001101110011101101011110010,
	240'b111010101011110011101000111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111111111111111111101001011101111100100,
	240'b101100101101000111111111111100011010010001111110011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111101101111000011110101001010111100011111111111110001110110011,
	240'b100100101110111011111110100110110100111001010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110110011110010100011100110100101101111100111101011111111010011011,
	240'b101010011111100111110011011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011000011101011111110100111010100111001101010101110101111111111110110000,
	240'b101101011111101111101101011000110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011111001111000010001100111001111001101001010001110100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011011001110110111011101111101101000010101010001110100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100101001111010111010100111100011011001001010100110100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100111011101001010000100101111110100001100110110011101111111110111100,
	240'b101101011111101111101101011001000101001101010011010100000101000101010010010100000100111101010001010100110101010001010101010101010101010101010101010101010101010001010111110101101011001101001100100100011110101001101000110011101111111110111100,
	240'b101101011111101111101101011001000100111101100010100101001010111110110000101010001001011101111110011000110101010001010000010101000101010101010101010101010101010101010001100111111111011011000111111011111011110101010110110100001111111110111100,
	240'b101101011111101111101101011000000111011011011010111111111111111111111111111111111111111111111001111001101011111110001001010110110101000001010100010101010101010101010100010110101010001011010010101100100110001101010100110100001111111110111100,
	240'b101101011111101111101010011101111110000011111111111111111111111111111111111111111111111111111111111111111111111111111100110101001000101101010110010100100101010101010101010101000101001001010111010100110101001001010110110100001111111110111100,
	240'b101101011111101111101001101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111000010011010110101000101010101010101010101010101010100010101010101010001010110110100001111111110111100,
	240'b101101011111100111110011111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011000001101010001010101000101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111100111111010111111001111111111111111111111111111111111111111111111111111111111111111111111111111111011101010111001111111101011111111111111111111001010001111010100010101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111100111111011111111011111111111111111111111111111111111111111111111111111111111111111111011101001010101100010010111111000001111011101111111111111111111110100100010110101000001010101010101010101010001010110110100001111111110111100,
	240'b101101011111100111111001111110001111111111111111111111111111111111111111111111111111111111111000100010110100111001001111010011100100111001110001111010101111111111111111111011110111100101010001010101010101010001010110110100001111111110111100,
	240'b101101011111100111110101111011011111111111111111111111111111111111111111111111111111111111001111010101010101001101111001100001000101011101001111101011011111111111111111111111111101101101100011010100110101010001010110110100001111111110111100,
	240'b101101011111101011101111110110111111111111111111111111111111111111111111111111111111111110101100010011100110010111100111111111000111110001001100100010111111111011111111111111111111111110110100010100110101010001010110110100001111111110111100,
	240'b101101011111101111101001110001001111111111111111111111111111111111111111111111111111111110101100010011100110010111100110111110100111101101001100100010111111111011111111111111111111111111110111011111010101000001010110110100001111111110111100,
	240'b101101011111101111101000101000101111111111111111111111111111111111111111111111111111111111010011010110100101001101110110100000010101011101010001101100011111111111111111111111111111111111111111110010010101011001010101110100001111111110111100,
	240'b101101011111101111101010100000011111001011111111111111111111111111111111111111111111111111100111011001110101001001010000010011110101001101011000110010111111111111111111111111111111111111111111111110010111110001010010110100001111111110111100,
	240'b101101011111101111101100011001111101000111111111111111111111111111111111111111111111101010001111010100100101001001011010010111010101001101010001011101011110110111111111111111111111111111111111111111111011100101010011110100001111111110111100,
	240'b101101011111101111101101010111111001111011111111111111111111111111111111111111111100110101010110010100011000001011010011110111001001101001010101010011111010110011111111111111111111111111111111111111111110100001100110110011101111111110111100,
	240'b101101011111101111101101011000010110100011101110111111111111111111111111111111111001110101001101011010001110100011111111111111111111101010000000010011000111110011111010111111111111111111111111111111111111110110001011110010111111111110111100,
	240'b101101011111101111101101011001000101000010110011111111111111111111111111111111111000100101001011100010011111111111111111111111111111111110101010010011010110110111110000111111111111111111111111111111111111111110110010110010111111111110111100,
	240'b101101011111101111101101011001000100111101101100111011011111111111111111111111111000111001001011100000011111110111111111111111111111111110100001010011000111000111110011111111111111111111111111111111111111111111010011110100111111111110111100,
	240'b101101011111101111101101011001000101001101010001101000001111111111111111111111111010110101001110010111001100110011111111111111111110010001101100010011011000100111111110111111111111111111111111111111111111111111101001110110111111111110111100,
	240'b101101011111101111101101011001000101001101010011010110101100111011111111111111111110001001100001010100000110010110100001101010010111000101010001010101001100010111111111111111111111111111111111111111111111111111110010111001111111111110111100,
	240'b101101011111101111101101011001000101001101010101010100010110111011100101111111111111111110110100010101010100111101010000010100000100111101010000100101011111101011111111111111111111111111111111111111111111111111110111111100001111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101000010000000111011101111111111111101101110010110111001010111010101110110010110100011111101101111111111111111111111111111111111111111111111111111111111111001111101011111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010000100001011110111011111111111111111110111111010010110011101110100011111111111111111111111111111111111111111111111111111111111111111111111111111010111101101111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010100010111110111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111010101111111110111100,
	240'b101101011111101111101101011001000101001101010101010101010101010101010101010101010101000001101100110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000110101011111111110111100,
	240'b101101011111101111101101011001000101001001010001010100100101000101010100010101010101010101010010010101111000111011011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001110110011001111111110111100,
	240'b101101011111101111101101011001000101001010001000101101101001100101011011010101000101010101010101010101000101000001011111100100001100101111110000111111101111111111111111111111111111111111111111111101101010001001010101110100001111111110111100,
	240'b101101011111101111101101011000001000101011110101111000101111011110101101010100110101010101010101010101010101010101010011010100000101011101101101100011111010101111000000110010111100111010111000011111100101001001010101110100001111111110111100,
	240'b101101011111101111101101011000111100111111000000010101101001110011101100011000110101001101010101010101010101010101010101010101010101010001010010010100000101000001010100010101110101100001010011010100010101010001010110110100001111111110111100,
	240'b101101011111101111101100011001001101011010110000010010001000100011110000011001100101001101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001010110110100001111111110111100,
	240'b101101011111101111101101011000001001111011110000101110011110010011000011010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111101111101101011000010110011111101110111100101111101110000111010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100001111111110111100,
	240'b101101011111101111101101011000000111100011101110100010101110000110011110010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100001111111110111101,
	240'b101011011111101011110001011001000110001111100010111001101111000101111111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110101001111111110110100,
	240'b100101011111000111111101100011010100101101111000101101101000110001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100111001110000111100001111111110011100,
	240'b101010001101100011111111111001101000100101100111011001100110011101101010011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010100111110011010010111111111110101010101011,
	240'b111001011011101111110001111111111111101111110001111100001111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100001111100011111111111110111011111011011101,
	240'b111100101110000010111101111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001101111111101000011110010,
	240'b111110011111101111100101101001011001011010101110101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001001110010011101110111101111110011111001,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule