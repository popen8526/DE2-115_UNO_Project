module blue_zero(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110101111001011100101101000001001101010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010000110011100111001011111111111101100,
	240'b111111001110001110110110110101101111010111110110111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101101111011011100010101111001110011011101111,
	240'b111101101011101011101010111111111111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111111111101101100000111011101,
	240'b110000001101011011111111111100001010011110001000100001101000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000010010000010100000111001100111100001111111111110101110110100,
	240'b100111101111010011111101100101000100111001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011100110100010010001011110010100110101110101111100011111111110101110,
	240'b101011001111111111101011011000110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011101101110011111110011111101101001111001010010110011001111111110101111,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011110000001101100101101111101011011110100101100100110000001111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101101010011101001001011101011110101101110101101111111111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101101010010101001101011101011110101001110101101111111111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101111010010101001100011101001110101001110101101111111111111110110000,
	240'b101100101111111111100010011000000101001101010011010100000101000101010001010011110101000001010001010100110101010101010101010101010101010101010101010101010101010001010110110011111011110001001110100001111110111001101110101111111111111110110001,
	240'b101100101111111111100010011000000100111101100011100100111010110110101101101000111001000101111001011000000101001101010000010101000101010101010101010101010101010101010001100101111111011111000110111010101100100001010110110000101111111110110001,
	240'b101100101111111111100010010111000111110111011110111111111111111111111111111111111111111111110111111000101011101010000110010110110101000001010100010101010101010101010100010110001001111011010110101110010110011101010010110000111111111110110001,
	240'b101100101111111111011111011110101110100011111111111111111111111111111111111111111111111111111111111111111111111111111100110101011000110101010111010100100101010101010101010101000101001001011000010101000101001001010100110000111111111110110001,
	240'b101100101111111111100000110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000100011011000101000001010101010101010101010101010100010101000101010001010100110000111111111110110001,
	240'b101100101111111111101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011000001101010001010101000101010101010101010101010101010001010100110000111111111110110001,
	240'b101100101111111111110011111110101111111111111111111111111111111111111111111111111111111111111111111111111111100111101000111001101111010011111111111111111111001110010011010100100101010001010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111110011111110011111111111111111111111111111111111111111111111111111111111111111110011011000000101100001010111100111010110111000111110101111111111110111100100110101000101010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111110001111110011111111111111111111111111111111111111111111111111111111111000000010110110100111101001110010011100100111101010011101000101111110011111111111101001000001001010000010101010101010001010100110000111111111110110000,
	240'b101100101111111111101101111100101111111111111111111111111111111111111111111111111110011101100111010011110101110010001010100100100110010101010001010101111100101011111111111111111110010001101010010100100101010001010100110000111111111110110000,
	240'b101100101111111111100111111000011111111111111111111111111111111111111111111111111011000001001111010110001011101111111110111111111101011001100110010011011000101111111110111111111111111111000000010101100101001101010100110000111111111110110000,
	240'b101100101111111111100000110010011111111111111111111111111111111111111111111111111000110101001100011111001111101111111111111111111111111110011110010011000110111011110100111111111111111111111011100010010100111101010100110000111111111110110001,
	240'b101100101111111111011101101010001111111111111111111111111111111111111111111111111000000101001010100011111111111111111111111111111111111110110011010011100110100011101100111111111111111111111111110101100101101001010011110000111111111110110001,
	240'b101100101111111111011110100000111111011111111111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111011000100101001111110000111111111110110001,
	240'b101100101111111111100001011001101101100011111111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111111100100001010100110000101111111110110001,
	240'b101100101111111111100010010110111010010011111111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111111111000101101101101111111111111110110001,
	240'b101100101111111111100010010111010110110011110001111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111111111111110010110101111011111111110110001,
	240'b101100101111111111100010011000000101000110110111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101100111111111111111111111111111111111111111110111111101111111111111110110000,
	240'b101100101111111111100010011000000101000001101110111011101111111111111111111111111000101101001011011111111111110011111111111111111111111110100010010011000110110111110011111111111111111111111111111111111111111111011100110010111111111110110000,
	240'b101100101111111111100010011000000101001101010001101000011111111111111111111111111010110101001111010110101100010111111111111111111101111101101010010011011000100011111101111111111111111111111111111111111111111111110000110101111111111110110000,
	240'b101100101111111111100010011000000101001101010011010110111100111111111111111111111110001101100100010100000110000010010111100111110110110001010001010101011100011011111111111111111111111111111111111111111111111111111000111000101111111110110000,
	240'b101100101111111111100010011000000101001101010101010100010110111011100101111111111111111110111001010110000100111101001111010011110100111101010001100110101111101111111111111111111111111111111111111111111111111111111010111010101111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101000001111111111011011111111111111111110000100111011001011101010110110110101110101100111110001111111111111111111111111111111111111111111111111111111111111011111011111111111110110001,
	240'b101100101111111111100010011000000101001101010101010101010101010101010000100000101110101111111111111111111111010111011110110110101110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111111111110110001,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010100010111011011011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111000111111111110110001,
	240'b101100101111111111100010011000000101001101010101010101000101010101010101010101010101000001100101101110011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011110010111111111110110001,
	240'b101100101111111111100010011000000101001001010001010101010101000101010100010101010101010101010010010101011000001111001101111110101111111111111111111111111111111111111111111111111111111111111111111111111111101010001110101111101111111110110001,
	240'b101100101111111111100010010111110101011110011011110010001010011001011101010100110101010101010101010101000101000001011001100000001011101011100101111110011111111111111111111111111111111111111111111100111001111101010011110000101111111110110001,
	240'b101100101111111111100010010111001001110111110110110100101111010010110010010100110101010101010101010101010101010101010100010100010101001101100010011111111001100010101110101110101011111010101001011110000101001001010011110000111111111110110000,
	240'b101100101111111111100001011000111101101010110010010011101001101111101010011000110101001101010101010101010101010101010101010101010101010001010011010100010101000001010010010100110101010001010001010100010101010001010100110000111111111110110000,
	240'b101100101111111111100001011010011110000010010110010010100111111111101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111100001011010011101111110010111010010111000000011101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111100001011010011110000010010110010010001000000011101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111100001011000011101001011000101011000101011000111100100010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110000101111111110110001,
	240'b101011011111111111101001010111101000011111110010111011011111011010011011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110010101111111110110000,
	240'b100111101111010111111100100011010100110001110111101000001000000001010010010100000101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100111001110000111011101111111110101110,
	240'b101111001101100111111111111010111001101001111000011101110111100001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011110111000110011011010111111111110110110110010,
	240'b111101001011100111101110111111111111111111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111111111111111110011100001111011010,
	240'b111110011110100010111101111000011111100011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111100111101001101111011101100111101000,
	240'b111101001111111111110010101001101000111010101101101100011011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001011010010000110101101111001111011111,
	240'b111110101111001011100101101000001001101010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010000110011100111001011111111111101100,
	240'b111111001110001110110110110101101111010111110110111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101101111011011100010101111001110011011101111,
	240'b111101101011101011101010111111111111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111111111101101100000111011101,
	240'b110000001101011011111111111100001010011110001000100001101000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000010010000010100000111001100111100001111111111110101110110100,
	240'b100111101111010011111101100101000100111001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011100110100010010001011110010100110101110101111100011111111110101110,
	240'b101011001111111111101011011000110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011101101110011111110011111101101001111001010010110011001111111110101111,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011110000001101100101101111101011011110100101100100110000001111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101101010011101001001011101011110101101110101101111111111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101101010010101001101011101011110101001110101101111111111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101111010010101001100011101001110101001110101101111111111111110110000,
	240'b101100101111111111100010011000000101001101010011010100000101000101010001010011110101000001010001010100110101010101010101010101010101010101010101010101010101010001010110110011111011110001001110100001111110111001101110101111111111111110110001,
	240'b101100101111111111100010011000000100111101100011100100111010110110101101101000111001000101111001011000000101001101010000010101000101010101010101010101010101010101010001100101111111011111000110111010101100100001010110110000101111111110110001,
	240'b101100101111111111100010010111000111110111011110111111111111111111111111111111111111111111110111111000101011101010000110010110110101000001010100010101010101010101010100010110001001111011010110101110010110011101010010110000111111111110110001,
	240'b101100101111111111011111011110101110100011111111111111111111111111111111111111111111111111111111111111111111111111111100110101011000110101010111010100100101010101010101010101000101001001011000010101000101001001010100110000111111111110110001,
	240'b101100101111111111100000110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000100011011000101000001010101010101010101010101010100010101000101010001010100110000111111111110110001,
	240'b101100101111111111101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011000001101010001010101000101010101010101010101010101010001010100110000111111111110110001,
	240'b101100101111111111110011111110101111111111111111111111111111111111111111111111111111111111111111111111111111100111101000111001101111010011111111111111111111001110010011010100100101010001010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111110011111110011111111111111111111111111111111111111111111111111111111111111111110011011000000101100001010111100111010110111000111110101111111111110111100100110101000101010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111110001111110011111111111111111111111111111111111111111111111111111111111000000010110110100111101001110010011100100111101010011101000101111110011111111111101001000001001010000010101010101010001010100110000111111111110110000,
	240'b101100101111111111101101111100101111111111111111111111111111111111111111111111111110011101100111010011110101110010001010100100100110010101010001010101111100101011111111111111111110010001101010010100100101010001010100110000111111111110110000,
	240'b101100101111111111100111111000011111111111111111111111111111111111111111111111111011000001001111010110001011101111111110111111111101011001100110010011011000101111111110111111111111111111000000010101100101001101010100110000111111111110110000,
	240'b101100101111111111100000110010011111111111111111111111111111111111111111111111111000110101001100011111001111101111111111111111111111111110011110010011000110111011110100111111111111111111111011100010010100111101010100110000111111111110110001,
	240'b101100101111111111011101101010001111111111111111111111111111111111111111111111111000000101001010100011111111111111111111111111111111111110110011010011100110100011101100111111111111111111111111110101100101101001010011110000111111111110110001,
	240'b101100101111111111011110100000111111011111111111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111011000100101001111110000111111111110110001,
	240'b101100101111111111100001011001101101100011111111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111111100100001010100110000101111111110110001,
	240'b101100101111111111100010010110111010010011111111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111111111000101101101101111111111111110110001,
	240'b101100101111111111100010010111010110110011110001111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101011111111111111111111111111111111111111111110010110101111011111111110110001,
	240'b101100101111111111100010011000000101000110110111111111111111111111111111111111111000000001001010100011111111111111111111111111111111111110110011010011100110100011101100111111111111111111111111111111111111111110111111101111111111111110110000,
	240'b101100101111111111100010011000000101000001101110111011101111111111111111111111111000101101001011011111111111110011111111111111111111111110100010010011000110110111110011111111111111111111111111111111111111111111011100110010111111111110110000,
	240'b101100101111111111100010011000000101001101010001101000011111111111111111111111111010110101001111010110101100010111111111111111111101111101101010010011011000100011111101111111111111111111111111111111111111111111110000110101111111111110110000,
	240'b101100101111111111100010011000000101001101010011010110111100111111111111111111111110001101100100010100000110000010010111100111110110110001010001010101011100011011111111111111111111111111111111111111111111111111111000111000101111111110110000,
	240'b101100101111111111100010011000000101001101010101010100010110111011100101111111111111111110111001010110000100111101001111010011110100111101010001100110101111101111111111111111111111111111111111111111111111111111111010111010101111111110110000,
	240'b101100101111111111100010011000000101001101010101010101010101000001111111111011011111111111111111110000100111011001011101010110110110101110101100111110001111111111111111111111111111111111111111111111111111111111111011111011111111111110110001,
	240'b101100101111111111100010011000000101001101010101010101010101010101010000100000101110101111111111111111111111010111011110110110101110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111111111110110001,
	240'b101100101111111111100010011000000101001101010101010101010101010101010101010100010111011011011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111000111111111110110001,
	240'b101100101111111111100010011000000101001101010101010101000101010101010101010101010101000001100101101110011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011110010111111111110110001,
	240'b101100101111111111100010011000000101001001010001010101010101000101010100010101010101010101010010010101011000001111001101111110101111111111111111111111111111111111111111111111111111111111111111111111111111101010001110101111101111111110110001,
	240'b101100101111111111100010010111110101011110011011110010001010011001011101010100110101010101010101010101000101000001011001100000001011101011100101111110011111111111111111111111111111111111111111111100111001111101010011110000101111111110110001,
	240'b101100101111111111100010010111001001110111110110110100101111010010110010010100110101010101010101010101010101010101010100010100010101001101100010011111111001100010101110101110101011111010101001011110000101001001010011110000111111111110110000,
	240'b101100101111111111100001011000111101101010110010010011101001101111101010011000110101001101010101010101010101010101010101010101010101010001010011010100010101000001010010010100110101010001010001010100010101010001010100110000111111111110110000,
	240'b101100101111111111100001011010011110000010010110010010100111111111101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111100001011010011101111110010111010010111000000011101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111100001011010011110000010010110010010001000000011101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110000111111111110110000,
	240'b101100101111111111100001011000011101001011000101011000101011000111100100010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110000101111111110110001,
	240'b101011011111111111101001010111101000011111110010111011011111011010011011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100110010101111111110110000,
	240'b100111101111010111111100100011010100110001110111101000001000000001010010010100000101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100111001110000111011101111111110101110,
	240'b101111001101100111111111111010111001101001111000011101110111100001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011110111000110011011010111111111110110110110010,
	240'b111101001011100111101110111111111111111111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111111111111111111110011100001111011010,
	240'b111110011110100010111101111000011111100011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111100111101001101111011101100111101000,
	240'b111101001111111111110010101001101000111010101101101100011011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001011010010000110101101111001111011111,
	240'b111110101111001011100101101000001001101010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001010000110011100111001011111111111101100,
	240'b111111001110001110110110110101101111010111110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101011111011011100010101111001110011011101111,
	240'b111101101011101011101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101100000111011101,
	240'b110000001101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010110100,
	240'b100111101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110,
	240'b101011001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101011011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b100111101111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110,
	240'b101111001101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110110010,
	240'b111101001011100111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100001111011010,
	240'b111110011110100010111101111000011111011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111100011101001101111011101100111101000,
	240'b111101001111111111110010101001101000111010101101101100011011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001011010010000110101101111001111011111,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule