module green_eight(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111011111111011111110001101010011001111010101010101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001110010100101111001111111001011110000,
	240'b111100001110101011000010110100101110110111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110101111001101101110111110100011110000,
	240'b111011001011110011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011011110111101110,
	240'b101111111101010011111111111100101010111010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001000010001101100100001011001011110110111111111100111110111110,
	240'b100100111111010111111100100101100100111001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011100110010110000001010111100100110110011111111111101111001010001101,
	240'b101001111111111011101001011000000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011010101101111111111011110100010101110001100111111011111111101010100011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111100101011110100110010000111100100111110001011110111010011111110010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100000101111001011010001111011110110110101011111111010011111110010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101001101111011011011111111101011001000001011110111010011111110010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111001011010001101010010101110001101001101100100111001111111110010110011,
	240'b101101101111111111100001010110110101010001010011010100000100111101001111010100000101000101010010010101000101010101010101010101010101010101010101010101010101001101100011111010011001010001001000101011001101100101100110111001111111110010110011,
	240'b101101101111111111100001010110110101000001100011100100111010101110101000100111101000100001110000010111000101000101010001010101000101010101010101010101010101010101010100101111001110110110111111111101001010010001011111111010001111110010110011,
	240'b101101101111111111100001010110000111110111011110111111111111111111111111111111111111110111110100110101111010110101110111010101100101000101010100010101010101010101010011011000111011100011011110101010110101101001100001111010011111110010110011,
	240'b101101101111111111011110011101111110100111111111111111111111111111111111111111111111111111111111111111111111111111110101110001110111101101010011010100110101010101010101010100110101001101010111010100100101001001100010111010011111110010110011,
	240'b101101101111111111011111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101111010111110101000101010101010101010101010101010100010101010101001101100010111010011111110010110011,
	240'b101101101111111011101111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110111000001010001010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111110111111001111111011111111111111111111111111111111111111111111111111111111111111111111111111111101111100110111001111111110111111111111111111110011001111010010100000101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111110111111010111111101111111111111111111111111111111111111111111111111111111111111111111000111000100101100011011001001000111011101000111111111111111111101000011110010101000001010101010101010101001101100010111010011111110010110011,
	240'b101101101111110111110111111110101111111111111111111111111111111111111111111111111111111111110000011110000100111001001111010011110100111010000000111101011111111111111111111000010110101001010010010101010101001101100010111010011111110010110011,
	240'b101101101111111011110001111100001111111111111111111111111111111111111111111111111111111110111001010100000101010110000010011111110101010001010010110001001111111111111111111111111100100101011001010101000101001101100010111010011111110010110011,
	240'b101101101111111111100111111000001111111111111111111111111111111111111111111111111111111110010111010011000111010111110110111100000110110001001100101000111111111111111111111111111111111110011101010100010101001101100010111010011111110010110011,
	240'b101101101111111111011111110010111111111111111111111111111111111111111111111111111111111110011000010011000111001011110001111010110110101001001100101001001111111111111111111111111111111111101011011010110101000001100010111010011111110010110011,
	240'b101101101111111111011100101010001111111111111111111111111111111111111111111111111111111111000010010101000101010001111000011101010101001101010111110011001111111111111111111111111111111111111111101100100101000001100010111010011111110010110011,
	240'b101101101111111111011101100001001111100111111111111111111111111111111111111111111111111111010011010110110101001101010000010100000101001101100000110111011111111111111111111111111111111111111111111011100110100101011111111010011111110010110011,
	240'b101101101111111111011111011001001101111011111111111111111111111111111111111111111111000001111000010100010101001001100000011000010101001001010001100000011111010111111111111111111111111111111111111111111001111101011101111010011111110010110011,
	240'b101101101111111111100001010101111010110011111111111111111111111111111111111111111011010101010000010101001001100111100000111000001001001101010010010100101100000011111111111111111111111111111111111111111101001101100110111001111111110010110011,
	240'b101101101111111111100001010110000111000111110100111111111111111111111111111111011000011101001100011110101111100011111111111111111111001101110001010011001001001011111111111111111111111111111111111111111111010010000001111001011111110010110011,
	240'b101101101111111111100001010110110101001010111101111111111111111111111111111110000111011001001100100111111111111111111111111111111111111110010011010010111000000111111011111111111111111111111111111111111111111110100010111000111111110010110011,
	240'b101101101111111111100001010110110101000001110011111100101111111111111111111110110111111001001100100100011111111111111111111111111111111110000110010010111000100011111101111111111111111111111111111111111111111111000110111001011111110010110011,
	240'b101101101111111111100001010110110101001101010001101001111111111111111111111111111001110101001101011000001101000111111111111111111100100001011100010011101010100011111111111111111111111111111111111111111111111111011110111010001111101110110011,
	240'b101101101111111111100001010110110101010001010011010111011101010011111111111111111101100001011100010100000110001110010110100101000110000001010000011000011110000011111111111111111111111111111111111111111111111111101011111100011111101010110011,
	240'b101101101111111111100001010110110101010001010101010100010111001011101001111111111111111010101101010101010100111001001110010011100100111001010111101101111111111111111111111111111111111111111111111111111111111111110010111101101111101010110011,
	240'b101101101111111111100001010110110101010001010101010101010101000010000011111100001111111111111101101111000111011001100001011000010111100111000011111111101111111111111111111111111111111111111111111111111111111111110110111110011111101010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010000100001111110110111111111111111111111010111100000111000011111011111111111111111111111111111111111111111111111111111111111111111111111111111110110111110011111101010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010100000111101011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111100001111101110110011,
	240'b101101101111111111100001010110110101010001010101010101000101010101010101010101010101000101100110101101111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111001011111110010110011,
	240'b101101101111111111100001010110110101001101010010010101010101001001010100010101010101010101010010010101001000000111001010111110011111111111111111111111111111111111111111111111111111111111111111111111111110001101110111111001101111110010110011,
	240'b101101101111111111100001010110100101110010101100110110001010110001011101010101000101010101010101010101000101000001011000011111111011100011100000111110101111111111111111111111111111111111111111110111100111100101011110111010011111110010110011,
	240'b101101101111111111100001010110011010110011110010110001101111001010101101010100100101010101010101010101010101010101010100010100010101001001100001011110001001001010100111101100011011000110010011011000100100111101100010111010011111110010110011,
	240'b101101101111111111011111011000011110010010100000010010001010000111100101010110110101010001010101010101010101010101010101010101010101010101010011010100010101000001010000010100000101000001010000010100110101001101100010111010011111110010110011,
	240'b101101101111111111011111011000001101111110101010010100001010101111100001010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111111111100001010110001001110111110100110110011111010110011110010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111111111100001010101110111011011110010110110001111001001110111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111111111100001010101101000100111101100100011011110110010001010010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101001111111111011101001010111010110010011011100111110011101110001100110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111011111111101010100011,
	240'b100100101111011011111100100100100100110001100110100010000110011001001101010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110100111110011100111111101111001010001100,
	240'b101110111101011111111111111100001010100010001010100010011000101110001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011011010110011110100111111111101000110111010,
	240'b111010111011101011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001011101111101100,
	240'b111110011110101110111011110101001110111111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111101111111001110110111010011101111111110111011111000,
	240'b111111111111110111100010101000001001101110110000101100111011001110110011101100111011001110110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110010101011111001101010101100111101011111111111111111,
	240'b111011111111011111110001101010011001111010101010101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001110010100101111001111111001011110000,
	240'b111100001110101011000010110100101110110111111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001110101111001101101110111110100011110000,
	240'b111011001011110011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011011110111101110,
	240'b101111111101010011111111111110011101011011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100011111000110110001111101100011111010111111111100111110111110,
	240'b100100111111010111111110110010101010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001101011001011000000101011111010011011001111111111111111001010001101,
	240'b101001111111110111110100101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101101011110111111111101111010001010111010110011111110001111100110100011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110010101111010011000111111110011011111010101110111101001111101010110011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110000011111100111101000111101111011011010101111111101001111101010110011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110100111111101111101111111110101100100010101110111101001111101010110011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100101101000110101001110111001110100110110001111101001111101010110011,
	240'b101101101111111011110000101011011010100110101001101010001010011110100111101001111010100010101000101010011010101010101010101010101010101010101010101010101010100110110001111101001100100110100011110101011110110010110010111101001111101010110011,
	240'b101101101111111011110000101011011010011110110001110010011101010111010011110011101100010010110111101011101010100010101000101010101010101010101010101010101010101010101001110111011111011011011111111110011101001010101111111101001111101010110011,
	240'b101101101111111011110000101010111011111011101111111111111111111111111111111111111111111011111010111010111101011010111011101010111010100010101010101010101010101010101001101100011101101111101111110101011010110110101111111101001111101010110011,
	240'b101101101111111011101111101110111111010011111111111111111111111111111111111111111111111111111111111111111111111111111010111000111011110110101001101010011010101010101010101010011010100110101011101010011010100010110000111101001111101010110011,
	240'b101101101111111011101111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010111101011111010100010101010101010101010101010101010101010101010100110110000111101001111101010110011,
	240'b101101101111110111110111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011011100010101000101010101010101010101010101010101010100110110000111101001111101010110011,
	240'b101101101111110111111100111111101111111111111111111111111111111111111111111111111111111111111111111111111111110111110010111100111111111011111111111111111111001010111100101010001010101010101010101010101010100110110000111101001111101010110011,
	240'b101101101111110111111100111111101111111111111111111111111111111111111111111111111111111111111111111100011100010010110001101100101100011111110100111111111111111111110100101111001010100010101010101010101010100110110000111101001111101010110011,
	240'b101101101111110111111011111111001111111111111111111111111111111111111111111111111111111111111000101111001010011010100111101001111010011010111111111110101111111111111111111100001011010010101000101010101010100110110000111101001111101010110011,
	240'b101101101111110111111000111101111111111111111111111111111111111111111111111111111111111111011100101010001010101011000001101111111010100110101000111000101111111111111111111111111110010010101100101010011010100110110000111101001111101010110011,
	240'b101101101111111011110011111100001111111111111111111111111111111111111111111111111111111111001011101001011011101011111011111110001011011010100110110100011111111111111111111111111111111111001110101010001010100110110000111101001111101010110011,
	240'b101101101111111011101111111001011111111111111111111111111111111111111111111111111111111111001100101001101011100011111000111101011011010010100110110100101111111111111111111111111111111111110101101101011010100010110000111101001111101010110011,
	240'b101101101111111011101110110101001111111111111111111111111111111111111111111111111111111111100000101010101010101010111011101110101010100110101011111001011111111111111111111111111111111111111111110110011010011110110000111101001111101010110011,
	240'b101101101111111011101110110000011111110011111111111111111111111111111111111111111111111111101001101011011010100110100111101001111010100110101111111011101111111111111111111111111111111111111111111101111011010010101111111101001111101010110011,
	240'b101101101111111011101111101100011110111011111111111111111111111111111111111111111111100010111100101010001010100110110000101100001010100110101000110000001111101011111111111111111111111111111111111111111100111110101110111101001111101010110011,
	240'b101101101111111011110000101010111101010111111111111111111111111111111111111111111101101010100111101010011100110011110000111011111100100110101001101010001101111111111111111111111111111111111111111111111110100110110010111101001111101010110011,
	240'b101101101111111011110000101010111011100011111001111111111111111111111111111111101100001110100110101111001111101111111111111111111111100110111000101001011100100011111111111111111111111111111111111111111111101010111111111100101111101010110011,
	240'b101101101111111011110000101011011010100111011110111111111111111111111111111111001011101010100101110011111111111111111111111111111111111111001001101001011100000011111101111111111111111111111111111111111111111111010001111100011111101010110011,
	240'b101101101111111011110000101011011010011110111001111110001111111111111111111111011011111010100101110010001111111111111111111111111111111111000010101001011100001111111110111111111111111111111111111111111111111111100010111100101111101010110011,
	240'b101101101111111011110000101011011010100110101000110100111111111111111111111111111100111010100110101011111110100011111111111111111110010010101101101001101101001111111111111111111111111111111111111111111111111111101111111101001111101010110011,
	240'b101101101111111011110000101011011010100110101001101011101110101011111111111111111110110010101101101010001011000111001011110010011010111110100111101100001111000011111111111111111111111111111111111111111111111111110101111110001111101010110011,
	240'b101101101111111011110000101011011010100110101010101010001011100111110100111111111111111111010110101010101010011110100111101001111010011110101011110110111111111111111111111111111111111111111111111111111111111111111000111110111111100110110011,
	240'b101101101111111011110000101011011010100110101010101010101010100011000001111101111111111111111110110111011011101110110000101100001011110011100001111111111111111111111111111111111111111111111111111111111111111111111010111111011111100110110011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101000110000111111011011111111111111111111101011110000111100001111101111111111111111111111111111111111111111111111111111111111111111111111111111111010111111001111100110110011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101010101010001011110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111110001111101010110011,
	240'b101101101111111011110000101011011010100110101010101010101010101010101010101010101010100010110011110110111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111100101111101010110011,
	240'b101101101111111011110000101011011010100010101000101010101010100010101001101010101010101010101001101010101100000011100101111111001111111111111111111111111111111111111111111111111111111111111111111111111111000110111011111100111111101010110011,
	240'b101101101111111011110000101011001010110111010101111010111101010110101110101010011010101010101010101010101010100010101100101111111101110011110000111111001111111111111111111111111111111111111111111011101011110010101111111101001111101010110011,
	240'b101101101111111011110000101011001101010111111000111000101111100011010110101010011010101010101010101010101010101010101001101010001010100010110000101110111100100111010011110110001101100011001001101100011010011110110000111101001111101010110011,
	240'b101101101111111011101111101100001111000111010000101000111101000011110010101011011010100110101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100110110000111101001111101010110011,
	240'b101101101111111011101111101100001110111111010100101001111101010111110000101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101010110011,
	240'b101101101111111011110000101010111100111011111010111011001111101011001111101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101010110011,
	240'b101101101111111011110000101010111011101111111001111011001111100110111011101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101010110011,
	240'b101101101111111011110000101010111100010011110101110001101111011011000101101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101010110011,
	240'b101001111111110111110100101011101011000111101110111111001110111010110010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110011111101111111100110100011,
	240'b100100101111010111111110110010011010010110110010110001001011001010100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011111001101111111111111001010001100,
	240'b101110111101011111111111111110001101001111000101110001001100010111000111110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101101011011111010111111111101000110111010,
	240'b111010111011101011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001011101111101100,
	240'b111110011110101110111011110101001110111111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001110110111010011101111111110111011111000,
	240'b111111111111110111100010101000001001101110110000101100111011001110110011101100111011001110110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110010101011111001101010101100111101011111111111111111,
	240'b111011111111011111110001101010011001111010101010101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001110010100101111001111111001011110000,
	240'b111100001110101011000010110100101110110111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110101111001101101110111110100011110000,
	240'b111011001011110011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011011110111101110,
	240'b101111111101010011111111111100101010111010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001000010001101100100001011001011110110111111111100111110111110,
	240'b100100111111010111111100100101100100111001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011100110010110000001010111100100110110011111111111101111001010001101,
	240'b101001111111111011101001011000000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011010101101111111111011110100010101110001100111111011111111101010100011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111100101011110100110010000111100100111110001011110111010011111110010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100000101111001011010001111011110110110101011111111010011111110010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101001101111011011011111111101011001000001011110111010011111110010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111001011010001101010010101110001101001101100100111001111111110010110011,
	240'b101101101111111111100001010110110101010001010011010100000100111101001111010100000101000101010010010101000101010101010101010101010101010101010101010101010101001101100011111010011001010001001000101011001101100101100110111001111111110010110011,
	240'b101101101111111111100001010110110101000001100011100100111010101110101000100111101000100001110000010111000101000101010001010101000101010101010101010101010101010101010100101111001110110110111111111101001010010001011111111010001111110010110011,
	240'b101101101111111111100001010110000111110111011110111111111111111111111111111111111111110111110100110101111010110101110111010101100101000101010100010101010101010101010011011000111011100011011110101010110101101001100001111010011111110010110011,
	240'b101101101111111111011110011101111110100111111111111111111111111111111111111111111111111111111111111111111111111111110101110001110111101101010011010100110101010101010101010100110101001101010111010100100101001001100010111010011111110010110011,
	240'b101101101111111111011111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101111010111110101000101010101010101010101010101010100010101010101001101100010111010011111110010110011,
	240'b101101101111111011101111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110111000001010001010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111110111111001111111011111111111111111111111111111111111111111111111111111111111111111111111111111101111100110111001111111110111111111111111111110011001111010010100000101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111110111111010111111101111111111111111111111111111111111111111111111111111111111111111111000111000100101100011011001001000111011101000111111111111111111101000011110010101000001010101010101010101001101100010111010011111110010110011,
	240'b101101101111110111110111111110101111111111111111111111111111111111111111111111111111111111110000011110000100111001001111010011110100111010000000111101011111111111111111111000010110101001010010010101010101001101100010111010011111110010110011,
	240'b101101101111111011110001111100001111111111111111111111111111111111111111111111111111111110111001010100000101010110000010011111110101010001010010110001001111111111111111111111111100100101011001010101000101001101100010111010011111110010110011,
	240'b101101101111111111100111111000001111111111111111111111111111111111111111111111111111111110010111010011000111010111110110111100000110110001001100101000111111111111111111111111111111111110011101010100010101001101100010111010011111110010110011,
	240'b101101101111111111011111110010111111111111111111111111111111111111111111111111111111111110011000010011000111001011110001111010110110101001001100101001001111111111111111111111111111111111101011011010110101000001100010111010011111110010110011,
	240'b101101101111111111011100101010001111111111111111111111111111111111111111111111111111111111000010010101000101010001111000011101010101001101010111110011001111111111111111111111111111111111111111101100100101000001100010111010011111110010110011,
	240'b101101101111111111011101100001001111100111111111111111111111111111111111111111111111111111010011010110110101001101010000010100000101001101100000110111011111111111111111111111111111111111111111111011100110100101011111111010011111110010110011,
	240'b101101101111111111011111011001001101111011111111111111111111111111111111111111111111000001111000010100010101001001100000011000010101001001010001100000011111010111111111111111111111111111111111111111111001111101011101111010011111110010110011,
	240'b101101101111111111100001010101111010110011111111111111111111111111111111111111111011010101010000010101001001100111100000111000001001001101010010010100101100000011111111111111111111111111111111111111111101001101100110111001111111110010110011,
	240'b101101101111111111100001010110000111000111110100111111111111111111111111111111011000011101001100011110101111100011111111111111111111001101110001010011001001001011111111111111111111111111111111111111111111010010000001111001011111110010110011,
	240'b101101101111111111100001010110110101001010111101111111111111111111111111111110000111011001001100100111111111111111111111111111111111111110010011010010111000000111111011111111111111111111111111111111111111111110100010111000111111110010110011,
	240'b101101101111111111100001010110110101000001110011111100101111111111111111111110110111111001001100100100011111111111111111111111111111111110000110010010111000100011111101111111111111111111111111111111111111111111000110111001011111110010110011,
	240'b101101101111111111100001010110110101001101010001101001111111111111111111111111111001110101001101011000001101000111111111111111111100100001011100010011101010100011111111111111111111111111111111111111111111111111011110111010001111101110110011,
	240'b101101101111111111100001010110110101010001010011010111011101010011111111111111111101100001011100010100000110001110010110100101000110000001010000011000011110000011111111111111111111111111111111111111111111111111101011111100011111101010110011,
	240'b101101101111111111100001010110110101010001010101010100010111001011101001111111111111111010101101010101010100111001001110010011100100111001010111101101111111111111111111111111111111111111111111111111111111111111110010111101101111101010110011,
	240'b101101101111111111100001010110110101010001010101010101010101000010000011111100001111111111111101101111000111011001100001011000010111100111000011111111101111111111111111111111111111111111111111111111111111111111110110111110011111101010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010000100001111110110111111111111111111111010111100000111000011111011111111111111111111111111111111111111111111111111111111111111111111111111111110110111110011111101010110011,
	240'b101101101111111111100001010110110101010001010101010101010101010101010101010100000111101011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111100001111101110110011,
	240'b101101101111111111100001010110110101010001010101010101000101010101010101010101010101000101100110101101111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111001011111110010110011,
	240'b101101101111111111100001010110110101001101010010010101010101001001010100010101010101010101010010010101001000000111001010111110011111111111111111111111111111111111111111111111111111111111111111111111111110001101110111111001101111110010110011,
	240'b101101101111111111100001010110100101110010101100110110001010110001011101010101000101010101010101010101000101000001011000011111111011100011100000111110101111111111111111111111111111111111111111110111100111100101011110111010011111110010110011,
	240'b101101101111111111100001010110011010110011110010110001101111001010101101010100100101010101010101010101010101010101010100010100010101001001100001011110001001001010100111101100011011000110010011011000100100111101100010111010011111110010110011,
	240'b101101101111111111011111011000011110010010100000010010001010000111100101010110110101010001010101010101010101010101010101010101010101010101010011010100010101000001010000010100000101000001010000010100110101001101100010111010011111110010110011,
	240'b101101101111111111011111011000001101111110101010010100001010101111100001010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111111111100001010110001001110111110100110110011111010110011110010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111111111100001010101110111011011110010110110001111001001110111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101101101111111111100001010101101000100111101100100011011110110010001010010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111010011111110010110011,
	240'b101001111111111011101001010111010110010011011100111110011101110001100110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111011111111101010100011,
	240'b100100101111011011111100100100100100110001100110100010000110011001001101010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110100111110011100111111101111001010001100,
	240'b101110111101011111111111111100001010100010001010100010011000101110001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011011010110011110100111111111101000110111010,
	240'b111010111011101011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001011101111101100,
	240'b111110011110101110111011110101001110111111111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111101111111001110110111010011101111111110111011111000,
	240'b111111111111110111100010101000001001101110110000101100111011001110110011101100111011001110110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110010101011111001101010101100111101011111111111111111,
};
assign data = picture[addr];
endmodule