module draw_card(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:49][29:0] picture = {
	30'b111111111111111111111111111111,
	30'b111111111111111111111111111111,
	30'b111111111111111111111111111111,
	30'b111000000000000000000000000111,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000010000000010000000011,
	30'b110000000010000000010000000011,
	30'b110000000010000001010000000011,
	30'b110000000010000000110000000011,
	30'b110000011111100000011110000011,
	30'b110000100010011000010000000011,
	30'b110000100010001000010000000011,
	30'b110000100010001000010000000011,
	30'b110001100010001011010000000011,
	30'b110001111111111000110000000011,
	30'b110000100010001000011100000011,
	30'b110000010010001000001011000011,
	30'b110000010010001000001001100011,
	30'b110000001010001000001000000011,
	30'b110000001100000000001000000011,
	30'b110000000011110000000110000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000010000000000011,
	30'b110000000011000010000000000011,
	30'b110000000000111100000000000011,
	30'b110000000000000100000000000011,
	30'b110000000000000100000000000011,
	30'b110000010000000010000000000011,
	30'b110000011111110010000000000011,
	30'b110000000000001111110000000011,
	30'b110000000000000001001110000011,
	30'b110000000000000010000000000011,
	30'b110000000000001110000000000011,
	30'b110000000000110010000000000011,
	30'b110000000011000010000000000011,
	30'b110000001100000010000000000011,
	30'b110000000000000010000000000011,
	30'b110000000000000010000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000011,
	30'b110000000000000000000000000111,
	30'b111000000000000000000000001111,
	30'b111111111111111111111111111111,
	30'b111111111111111111111111111111
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = {8{picture[(y_cnt - y_pin)][(x_cnt - x_pin)]}};
        g_data = {8{picture[(y_cnt - y_pin)][(x_cnt - x_pin)]}};
        b_data = {8{picture[(y_cnt - y_pin)][(x_cnt - x_pin)]}};
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule