module blue_two(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111111001111001111011101100111011010011011000001110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000011101111101001111110110011111110001111111111111011,
	240'b111111101110100110111011110010011110001111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001110000011000011110100001111111011111100,
	240'b111110111011110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001101001111111101,
	240'b110011011101001111111111111101011011110010100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011001111010011100101000111100101111111101111111101100011111001100,
	240'b101001001111011011111100100110000101000001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010011110110011101111001010110010101010010111100111111111110000110100000,
	240'b101011001111111111100100010111110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100011011110110011110101110100100110001001111000111110111111001010110001,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111000111011110110000101111010101010111101101100111101001111010110111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110010111011110111011101001000100110011010011101110000111100111111010110111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101011100001010111010100100101001101110001111101001111010110111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000101110110111000011011001010100110101110001111101001111010110111000,
	240'b101100011111111111010111010110100101010001010011010100000101000001010000010011110101000001010010010101000101010101010101010101010101010101010101010101010101010101011001011001000111110111100000110111110111100001101111111101001111010110111000,
	240'b101100011111111111010111010110100101000001100010100010101010000010011101100100101000000001101010010101110101000001010010010101000101010101010101010101010101001001110000111000111011001110111111111111111100100001110000111100111111010110111000,
	240'b101100011111111111010111010101110111111111011100111111111111111111111111111111111111101011101101110011111010001101110000010100110101000101010101010101010101001001101101110110101110001111100000111000001011000001110001111100111111010110111000,
	240'b101100011111111111010011011110011110101111111111111111111111111111111111111111111111111111111111111111111111111111110000101110010111000101010001010101000101010101010110010111010101111001011110010111100101100001110001111101001111010110111000,
	240'b101100011111111111010110110001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110100000010110010101001001010101010100110101001101010011010100110101000101110001111101001111010110111000,
	240'b101100011111111111100110111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001010110010101010001010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111110000111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111010011111001111111111111111111101100101101110010100010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111110001111110011111111111111111111111111111111111111111111111111111111111111111111001001001010101101000011000000111000010101100111101011111111111011101011011000101000101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111101101111110001111111111111111111111111111111111111111111111111111111111011111011011100100111001001110010011010100111001010000100011001111011011111111110101000110000101010011010101010101001001110001111101001111010110111000,
	240'b101100011111111111101000111101011111111111111111111111111111111111111111111111111111101010000110010011100101010101111111100101010110111101010001010100001011001011111111111111111011100001010100010101000101001001110001111101001111010110111000,
	240'b101100011111111111100000111010001111111111111111111111111111111111111111111111111101100101011010010100011001101111111000111111111110100001111000010011100111010111110110111111111111101110001101010100000101001001110001111101001111010110111000,
	240'b101100011111111111011000110100011111111111111111111111111111111111111111111111111011101001001111011000101110011011111111111111111111111110111100010011000101101011100011111111111111111111100000011000100100111101110001111101001111010110111000,
	240'b101100011111111111010010101100001111111111111111111111111111111111111111111111111011001001001100011010011111000011111111111111111111111111011011011111001000000011100011111111111111111111111111101000010100110101110001111101001111010110111000,
	240'b101100011111111111010010100010101111110011111111111111111111111111111111111111111100010101010010010101111100110111111111111111111111111111111101111110011111100111111101111111111111111111111111111000100101110101101111111101001111010110111000,
	240'b101100011111111111010101011001111110010011111111111111111111111111111111111111111110101101101000010011100111101011101000111111111111111111111111111111111111111111111111111111111111111111111111111111101000110101101011111101001111010110111000,
	240'b101100011111111111010111010101111011001111111111111111111111111111111111111111111111111110110101010101010100111101110011110101101111111111111111111111111111111111111111111111111111111111111111111111111100000101101111111100111111010110111000,
	240'b101100011111111111010111010101100111011011110111111111111111111111111111111111111111111111111101101011010101011101001110011000011011011111111011111111111111111111111111111111111111111111111111111111111110100010000011111100101111010110111000,
	240'b101100011111111111010111010110100101001111000010111111111111111111111111111111111111111111111111111111111011101001011101010011100101010010001111111010101111111111111111111111111111111111111111111111111111101010100001111011111111010110111000,
	240'b101100011111111111010111010110100101000001110110111101001111111111111111111111111111111111111111111111111111111111001110011011110100111101010000011100101100111011111110111111111111111111111111111111111111111111000001111011111111010110111000,
	240'b101100011111111111010111010110100101010001010010101010111111111111111111111111111100011110000010100110011111101011111111111010001000101001010101010011110110001111100011111111111111111111111111111111111111111111011011111100011111010110111000,
	240'b101100011111111111010111010110100101010001010011010111111101011111111111111111111010110101001000010110011001000110010110100110011000110001011011010100110101101011011001111111111111111111111111111111111111111111101101111100111111010010111000,
	240'b101100011111111111010111010110100101010001010101010100010111001111101010111111111010111001001101010100100100111001001110010011100101000001010011010100100101100111011001111111111111111111111111111111111111111111110010111101101111010010111000,
	240'b101100011111111111010111010110100101010001010101010101010101000010000011111100111011101101100000011001010110010101100101011001010110010101100101011001000110101111011110111111111111111111111111111111111111111111110100111101111111010010111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010000100001101110000111101001111001101110011011100110111001101110011011100110111001101110011111111010111111111111111111111111111111111111111111110100111101111111010010111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010100000111100011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110111100101111010110111000,
	240'b101100011111111111010111010110100101001001010011010100110101001101010011010101010101000101100011101101001111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010111011111111010110111000,
	240'b101100011111111111010111010111000110000001100011011000110110001101100000010101010101010101010010010101000111110011000100111101001111111111111111111111111111111111111111111111111111111111111111111111111100100101111000111100111111010110111000,
	240'b101100011111111111010101011010011100111111100010111000111110011011000110010110100101010001010101010101000101000101010101011101101010101111010110111100001111110111111111111111111111111111111010110001100110001101101110111101001111010110111000,
	240'b101100011111111111010100011010111110110011110100101010111100000011001110010110100101010001010101010101010101010101010100010100010101000101011010011011101000000110010101100111101001110001111110010110010100111101110001111101001111010110111000,
	240'b101100011111111111010111010110101000111111101011110011000110110101011110010101100101010101010101010101010101010101010101010101010101010101010100010100100101000101010000010100000101000001010001010101000101001001110001111101001111010110111000,
	240'b101100011111111111010111010110010100111001110100110110101101110101101100010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111010111010110110101011001010000011000011101011111000001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111010101011001111100001101111100010001101010000111011101010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111010110010111101101011111001111100000111101110111000001010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110000111101001111010110111000,
	240'b101011001111111111100100010111000111101111100100111101101101101101110000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111101111011111110111111001010110001,
	240'b101001001111010111111101100110110100111101100000011101010101110001001101010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101100110111110111111111110000010100000,
	240'b110100001101000111111111111110001011111110100101101001001010011010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001100111011111110111111101100011111001111,
	240'b111111001011110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101101010111111101,
	240'b111101011111010111001000110010011101011111011011110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110111101010111000000110010011111001011110101,
	240'b111100101111111111101010101000011001111010111001101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101101011001011010101001111001111111000011110011,
	240'b111111001111001111011101100111011010011011000001110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000011101111101001111110110011111110001111111111111011,
	240'b111111101110100110111011110010011110001111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001110000011000011110100001111111011111100,
	240'b111110111011110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001101001111111101,
	240'b110011011101001111111111111101011011110010100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011001111010011100101000111100101111111101111111101100011111001100,
	240'b101001001111011011111100100110000101000001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010011110110011101111001010110010101010010111100111111111110000110100000,
	240'b101011001111111111100100010111110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100011011110110011110101110100100110001001111000111110111111001010110001,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111000111011110110000101111010101010111101101100111101001111010110111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110010111011110111011101001000100110011010011101110000111100111111010110111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101011100001010111010100100101001101110001111101001111010110111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000101110110111000011011001010100110101110001111101001111010110111000,
	240'b101100011111111111010111010110100101010001010011010100000101000001010000010011110101000001010010010101000101010101010101010101010101010101010101010101010101010101011001011001000111110111100000110111110111100001101111111101001111010110111000,
	240'b101100011111111111010111010110100101000001100010100010101010000010011101100100101000000001101010010101110101000001010010010101000101010101010101010101010101001001110000111000111011001110111111111111111100100001110000111100111111010110111000,
	240'b101100011111111111010111010101110111111111011100111111111111111111111111111111111111101011101101110011111010001101110000010100110101000101010101010101010101001001101101110110101110001111100000111000001011000001110001111100111111010110111000,
	240'b101100011111111111010011011110011110101111111111111111111111111111111111111111111111111111111111111111111111111111110000101110010111000101010001010101000101010101010110010111010101111001011110010111100101100001110001111101001111010110111000,
	240'b101100011111111111010110110001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110100000010110010101001001010101010100110101001101010011010100110101000101110001111101001111010110111000,
	240'b101100011111111111100110111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001010110010101010001010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111110000111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111010011111001111111111111111111101100101101110010100010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111110001111110011111111111111111111111111111111111111111111111111111111111111111111001001001010101101000011000000111000010101100111101011111111111011101011011000101000101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111101101111110001111111111111111111111111111111111111111111111111111111111011111011011100100111001001110010011010100111001010000100011001111011011111111110101000110000101010011010101010101001001110001111101001111010110111000,
	240'b101100011111111111101000111101011111111111111111111111111111111111111111111111111111101010000110010011100101010101111111100101010110111101010001010100001011001011111111111111111011100001010100010101000101001001110001111101001111010110111000,
	240'b101100011111111111100000111010001111111111111111111111111111111111111111111111111101100101011010010100011001101111111000111111111110100001111000010011100111010111110110111111111111101110001101010100000101001001110001111101001111010110111000,
	240'b101100011111111111011000110100011111111111111111111111111111111111111111111111111011101001001111011000101110011011111111111111111111111110111100010011000101101011100011111111111111111111100000011000100100111101110001111101001111010110111000,
	240'b101100011111111111010010101100001111111111111111111111111111111111111111111111111011001001001100011010011111000011111111111111111111111111011011011111001000000011100011111111111111111111111111101000010100110101110001111101001111010110111000,
	240'b101100011111111111010010100010101111110011111111111111111111111111111111111111111100010101010010010101111100110111111111111111111111111111111101111110011111100111111101111111111111111111111111111000100101110101101111111101001111010110111000,
	240'b101100011111111111010101011001111110010011111111111111111111111111111111111111111110101101101000010011100111101011101000111111111111111111111111111111111111111111111111111111111111111111111111111111101000110101101011111101001111010110111000,
	240'b101100011111111111010111010101111011001111111111111111111111111111111111111111111111111110110101010101010100111101110011110101101111111111111111111111111111111111111111111111111111111111111111111111111100000101101111111100111111010110111000,
	240'b101100011111111111010111010101100111011011110111111111111111111111111111111111111111111111111101101011010101011101001110011000011011011111111011111111111111111111111111111111111111111111111111111111111110100010000011111100101111010110111000,
	240'b101100011111111111010111010110100101001111000010111111111111111111111111111111111111111111111111111111111011101001011101010011100101010010001111111010101111111111111111111111111111111111111111111111111111101010100001111011111111010110111000,
	240'b101100011111111111010111010110100101000001110110111101001111111111111111111111111111111111111111111111111111111111001110011011110100111101010000011100101100111011111110111111111111111111111111111111111111111111000001111011111111010110111000,
	240'b101100011111111111010111010110100101010001010010101010111111111111111111111111111100011110000010100110011111101011111111111010001000101001010101010011110110001111100011111111111111111111111111111111111111111111011011111100011111010110111000,
	240'b101100011111111111010111010110100101010001010011010111111101011111111111111111111010110101001000010110011001000110010110100110011000110001011011010100110101101011011001111111111111111111111111111111111111111111101101111100111111010010111000,
	240'b101100011111111111010111010110100101010001010101010100010111001111101010111111111010111001001101010100100100111001001110010011100101000001010011010100100101100111011001111111111111111111111111111111111111111111110010111101101111010010111000,
	240'b101100011111111111010111010110100101010001010101010101010101000010000011111100111011101101100000011001010110010101100101011001010110010101100101011001000110101111011110111111111111111111111111111111111111111111110100111101111111010010111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010000100001101110000111101001111001101110011011100110111001101110011011100110111001101110011111111010111111111111111111111111111111111111111111110100111101111111010010111000,
	240'b101100011111111111010111010110100101010001010101010101010101010101010101010100000111100011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110111100101111010110111000,
	240'b101100011111111111010111010110100101001001010011010100110101001101010011010101010101000101100011101101001111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110010111011111111010110111000,
	240'b101100011111111111010111010111000110000001100011011000110110001101100000010101010101010101010010010101000111110011000100111101001111111111111111111111111111111111111111111111111111111111111111111111111100100101111000111100111111010110111000,
	240'b101100011111111111010101011010011100111111100010111000111110011011000110010110100101010001010101010101000101000101010101011101101010101111010110111100001111110111111111111111111111111111111010110001100110001101101110111101001111010110111000,
	240'b101100011111111111010100011010111110110011110100101010111100000011001110010110100101010001010101010101010101010101010100010100010101000101011010011011101000000110010101100111101001110001111110010110010100111101110001111101001111010110111000,
	240'b101100011111111111010111010110101000111111101011110011000110110101011110010101100101010101010101010101010101010101010101010101010101010101010100010100100101000101010000010100000101000001010001010101000101001001110001111101001111010110111000,
	240'b101100011111111111010111010110010100111001110100110110101101110101101100010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111010111010110110101011001010000011000011101011111000001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111010101011001111100001101111100010001101010000111011101010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110001111101001111010110111000,
	240'b101100011111111111010110010111101101011111001111100000111101110111000001010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001110000111101001111010110111000,
	240'b101011001111111111100100010111000111101111100100111101101101101101110000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111101111011111110111111001010110001,
	240'b101001001111010111111101100110110100111101100000011101010101110001001101010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101100110111110111111111110000010100000,
	240'b110100001101000111111111111110001011111110100101101001001010011010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001100111011111110111111101100011111001111,
	240'b111111001011110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101101010111111101,
	240'b111101011111010111001000110010011101011111011011110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110111101010111000000110010011111001011110101,
	240'b111100101111111111101010101000011001111010111001101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101101011001011010101001111001111111000011110011,
	240'b111111001111001111011101100111011010011011000001110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000011101111101001111110110011111110001111111111111011,
	240'b111111101110100110111011110010011110001011100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001110000011000011110100001111111011111100,
	240'b111110111011110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100001101001111111101,
	240'b110011011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011111001100,
	240'b101001001111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110100000,
	240'b101011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110110001,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111000,
	240'b101011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110110001,
	240'b101001001111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010100000,
	240'b110100001101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011111001111,
	240'b111111001011110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011101101010111111101,
	240'b111101011111010111001000110010011101011111011011110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110111101010111000000110010011111001011110101,
	240'b111100101111111111101010101000011001111010111001101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101101011001011010101001111001111111000011110011,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule