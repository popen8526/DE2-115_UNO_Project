module red_three(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
    240'b111100011111101011011100101101101011000010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011000010110101110110011111000111101110,
    240'b111101101101100111000011111011011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011101001101111001101010011110010,
    240'b110110111100010011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011011110011011111,
    240'b101100101111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110110001,
    240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100101,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010,
    240'b101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001,
    240'b101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010,
    240'b101100011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110101010,
    240'b110011011101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011011010011,
    240'b111100111100100111010101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110011001100010011110001,
    240'b111110001111011011000101101011101011101111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100110110000110011001111011011110110,
    240'b111100011111101011011101101101101011000110110011101100101011001010110010101100101011001110110011101100111011001110110011101100111011001010110010101100101011001010110011101100111011001110110011101100111011000010110101110110101111000111101110,
    240'b111101101101100111000011111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001101111001101010011110010,
    240'b110110111100010011111100111111111111101111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100111111110111111111111110011011110011011111,
    240'b101100101111000011111111110100101000010001110010011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100100110111101101110011011111000101011011101111111111110011110110001,
    240'b101101011111111111101011011010110100111001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100000111001110100010011110010100110001111000111101001111111010100101,
    240'b101110011111111111000110010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011010101110010011110000111100010111011001010100110110001111111110110111,
    240'b101110011111111110111110010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001111111000010000010101001110111100101010100110100001111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011101001111010011011100011101000100111001010111110100011111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101001011111010011001000011100100100111001010111110100011111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011111000011010101001001111010110000110100001011010110100011111111110111010,
    240'b101110011111111110111111010100110101010001010010010100000101001101010010010100000101000001010001010100110101010101010101010101010101010101010101010101010101010001011011111000011010100101001110100101101101100001100010110011111111111110111010,
    240'b101110011111111110111111010100100101001001110011101001011011011010110100101010111001011101111100011000010101001101010001010101000101010101010101010101010101010101010010101001111111011011001011111101001011011101010110110100011111111110111010,
    240'b101110011111111110111110010100101001101011101111111111111111111111111111111111111111111111111000111000101011100110000010010110000101000101010100010101010101010101010100010111001010001111001111101010110101111101010101110100011111111110111010,
    240'b101110011111111110111011100010111111101011111111111111111111111111111111111111111111111111111111111111111111111111111001110011011000001101010100010100100101010101010101010101000101001001010110010100100101001001010111110100011111111110111010,
    240'b101110011111111111000111110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111001011001010101000101010101010101010101010101010100010101010101010001010111110100011111111110111010,
    240'b101110011111111111100000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010111100101010000010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111101101111111001111111111111111111111111111111111111111111111111111111111111111111111111111101011100111111010011111110111111111111111111110101110000100010100010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111101110111111001111111111111111111111111111111111111111111111111111111111111111110111111000011001011111011000011000111111101000111111111111111111101111100000010101000001010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111101010111110111111111111111111111111111111111111111111111111111111111111101100011101000100111001001111010011110100111010000000111101001111111111111111111010000111000101010001010101010101010001010111110100011111111110111010,
    240'b101110011111111111100011111110011111111111111111111111111111111111111111111111111111111110101111010011110101011001111111011110100101001001010000110000001111111111111111111111111101001001011110010100110101010001010111110100011111111110111010,
    240'b101110011111111111010111111100101111111111111111111111111111111111111111111111111111111110001011010010110111011111111000111011000111011001011100101001101111111111111111111111111111111110101001010100100101010001010111110100011111111110111010,
    240'b101110011111111111001011111000011111111111111111111111111111111111111111111111111111111110001011010010110111100011111000111111111111010011101100111101001111111111111111111111111111111111110011011101010101000001010111110100011111111110111010,
    240'b101110011111111110111101110001011111111111111111111111111111111111111111111111111111111110110000010100010101011010000010100101011101010011111111111111111111111111111111111111111111111111111111110000000101001101010111110100011111111110111010,
    240'b101110011111111110111010100111101111111111111111111111111111111111111111111111111111111111001110010110010101001101001111010010101011010011111111111111111111111111111111111111111111111111111111111101100111010101010011110100011111111110111010,
    240'b101110011111111110111011011100111111011011111111111111111111111111111111111111111111000001111001010100100101001001011001010110011011101011111111111111111111111111111111111111111111111111111111111111111011000101010011110100011111111110111010,
    240'b101110011111111110111110010101111101001011111111111111111111111111111111111111111011000001010000010100111000110111010010110111101111000111111111111111111111111111111111111111111111111111111111111111111110001101100011110011111111111110111010,
    240'b101110011111111110111111010011101001010111111111111111111111111111111111111111000111110001001101011110011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110000110110011001111111110111010,
    240'b101110011111111110111111010100010110000111100001111111111111111111111111111100010110101101001101101001011111111111111111111111111111111111101101110111101110011011111110111111111111111111111111111111111111111110101101110011001111111110111010,
    240'b101110011111111110111111010100110100111110010111111111101111111111111111111100110110111001001100101000001111111111111111111111111111111110010100010101101000001111111101111111111111111111111111111111111111111111001111110100011111111110111010,
    240'b101110011111111110111111010100110101001101011100110100001111111111111111111111011000010101001101011011101110100011111111111111111101110101100011010010111001011011111111111111111111111111111111111111111111111111100101110111011111111110111010,
    240'b101110011111111110111111010100110101010001010001011101111111000111111111111111111011111001010010010100100111100010110110101100100111000001010001010101111100111011111111111111111111111111111111111111111111111111110100111010001111111110111010,
    240'b101110011111111110111111010100110101010001010101010100011001011111111011111111111111100010001100010011110101000001010010010100010101000001010000100110101111110011111111111111111111111111111111111111111111111111111100111011101111111110111010,
    240'b101110011111111110111111010100110101010001010101010101000101010010101100111111101111111111110001100101100101111001010010010100110110000110100001111101101111111111111111111111111111111111111111111111111111111111111100111100011111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101001101010111101100001111111011111111111111101101110110111111110000011110000111111111111111111111111111111111111111111111111111111111111111111111111111111100111100101111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010011010101101010010011111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011001111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101000101001110001011111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110110011111111110111010,
    240'b101110011111111110111111010100110101001101010001010100010101001001010101010101010101010001010000011010001011000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010111110011011111111110111010,
    240'b101110011111111110111111010100100101011110001000100111110111010101010011010101010101010101010101010100100101001001110011101011111110001111111101111111111111111111111111111111111111111111111111111111001011000001011001110100001111111110111010,
    240'b101110011111111110111111010100101010100011111001111100011110111001111101010100010101010101010101010101010101010101010010010100100110001110000011101010011100010111010110110111101110000011001011100011100101010101010110110100011111111110111010,
    240'b101110011111111110111101011001101110100110100011011001101101001011000110010101000101010001010101010101010101010101010101010101010101001101010001010100000101001101011100011000000110000101010111010100010101001101010111110100011111111110111010,
    240'b101110011111111110111110010111101000010001011011010010001011000011010101010101110101010001010101010101010101010101010101010101010101010101010101010101010101010001010100010100110101001101010100010101010101010001010111110100011111111110111010,
    240'b101110011111111110111111010100100100111001101101101000001110101110101011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111110111111010100110100111010010000111110111110111001101011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111110111111010100010110111110000101100011101111001001110011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111000001010011101001001011101111110100011110101101101010010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110101001111111110111001,
    240'b101101111111111111011110010111000101100010101110110101001000110001010010010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101000001100111111010111111111110101010,
    240'b101100011111100011111110101100010110000101011000010111010101100001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100110011110111111111111111111000110101010,
    240'b110011011101000011111111111111111110010111011001110110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110011110100011111111111111111100011011010011,
    240'b111100111100100111010101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110011001100010011110001,
    240'b111110001111011011000101101011101011101111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100110110000110011001111011011110110,
    240'b111100011111101011011100101101101011000010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011000010110101110110011111000111101110,
    240'b111101101101100111000011111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001101111001101010011110010,
    240'b110110111100010011111100111111111111101111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100111111110111111111111110011011110011011111,
    240'b101100101111000011111111110100101000010001110010011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100100110111101101110011011111000101011011101111111111110011110110001,
    240'b101101011111111111101011011010110100111001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100000111001110100010011110010100110001111000111101001111111010100101,
    240'b101110011111111111000110010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011010101110010011110000111100010111011001010100110110001111111110110111,
    240'b101110011111111110111110010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001111111000010000010101001110111100101010100110100001111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011101001111010011011100011101000100111001010111110100011111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101001011111010011001000011100100100111001010111110100011111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011111000011010101001001111010110000110100001011010110100011111111110111010,
    240'b101110011111111110111111010100110101010001010010010100000101001101010010010100000101000001010001010100110101010101010101010101010101010101010101010101010101010001011011111000011010100101001110100101101101100001100010110011111111111110111010,
    240'b101110011111111110111111010100100101001001110011101001011011011010110100101010111001011101111100011000010101001101010001010101000101010101010101010101010101010101010010101001111111011011001011111101001011011101010110110100011111111110111010,
    240'b101110011111111110111110010100101001101011101111111111111111111111111111111111111111111111111000111000101011100110000010010110000101000101010100010101010101010101010100010111001010001111001111101010110101111101010101110100011111111110111010,
    240'b101110011111111110111011100010111111101011111111111111111111111111111111111111111111111111111111111111111111111111111001110011011000001101010100010100100101010101010101010101000101001001010110010100100101001001010111110100011111111110111010,
    240'b101110011111111111000111110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111001011001010101000101010101010101010101010101010100010101010101010001010111110100011111111110111010,
    240'b101110011111111111100000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010111100101010000010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111101101111111001111111111111111111111111111111111111111111111111111111111111111111111111111101011100111111010011111110111111111111111111110101110000100010100010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111101110111111001111111111111111111111111111111111111111111111111111111111111111110111111000011001011111011000011000111111101000111111111111111111101111100000010101000001010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111101010111110111111111111111111111111111111111111111111111111111111111111101100011101000100111001001111010011110100111010000000111101001111111111111111111010000111000101010001010101010101010001010111110100011111111110111010,
    240'b101110011111111111100011111110011111111111111111111111111111111111111111111111111111111110101111010011110101011001111111011110100101001001010000110000001111111111111111111111111101001001011110010100110101010001010111110100011111111110111010,
    240'b101110011111111111010111111100101111111111111111111111111111111111111111111111111111111110001011010010110111011111111000111011000111011001011100101001101111111111111111111111111111111110101001010100100101010001010111110100011111111110111010,
    240'b101110011111111111001011111000011111111111111111111111111111111111111111111111111111111110001011010010110111100011111000111111111111010011101100111101001111111111111111111111111111111111110011011101010101000001010111110100011111111110111010,
    240'b101110011111111110111101110001011111111111111111111111111111111111111111111111111111111110110000010100010101011010000010100101011101010011111111111111111111111111111111111111111111111111111111110000000101001101010111110100011111111110111010,
    240'b101110011111111110111010100111101111111111111111111111111111111111111111111111111111111111001110010110010101001101001111010010101011010011111111111111111111111111111111111111111111111111111111111101100111010101010011110100011111111110111010,
    240'b101110011111111110111011011100111111011011111111111111111111111111111111111111111111000001111001010100100101001001011001010110011011101011111111111111111111111111111111111111111111111111111111111111111011000101010011110100011111111110111010,
    240'b101110011111111110111110010101111101001011111111111111111111111111111111111111111011000001010000010100111000110111010010110111101111000111111111111111111111111111111111111111111111111111111111111111111110001101100011110011111111111110111010,
    240'b101110011111111110111111010011101001010111111111111111111111111111111111111111000111110001001101011110011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110000110110011001111111110111010,
    240'b101110011111111110111111010100010110000111100001111111111111111111111111111100010110101101001101101001011111111111111111111111111111111111101101110111101110011011111110111111111111111111111111111111111111111110101101110011001111111110111010,
    240'b101110011111111110111111010100110100111110010111111111101111111111111111111100110110111001001100101000001111111111111111111111111111111110010100010101101000001111111101111111111111111111111111111111111111111111001111110100011111111110111010,
    240'b101110011111111110111111010100110101001101011100110100001111111111111111111111011000010101001101011011101110100011111111111111111101110101100011010010111001011011111111111111111111111111111111111111111111111111100101110111011111111110111010,
    240'b101110011111111110111111010100110101010001010001011101111111000111111111111111111011111001010010010100100111100010110110101100100111000001010001010101111100111011111111111111111111111111111111111111111111111111110100111010001111111110111010,
    240'b101110011111111110111111010100110101010001010101010100011001011111111011111111111111100010001100010011110101000001010010010100010101000001010000100110101111110011111111111111111111111111111111111111111111111111111100111011101111111110111010,
    240'b101110011111111110111111010100110101010001010101010101000101010010101100111111101111111111110001100101100101111001010010010100110110000110100001111101101111111111111111111111111111111111111111111111111111111111111100111100011111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101001101010111101100001111111011111111111111101101110110111111110000011110000111111111111111111111111111111111111111111111111111111111111111111111111111111100111100101111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010011010101101010010011111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011001111111110111010,
    240'b101110011111111110111111010100110101010001010101010101010101010101010101010101000101001110001011111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110110011111111110111010,
    240'b101110011111111110111111010100110101001101010001010100010101001001010101010101010101010001010000011010001011000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010111110011011111111110111010,
    240'b101110011111111110111111010100100101011110001000100111110111010101010011010101010101010101010101010100100101001001110011101011111110001111111101111111111111111111111111111111111111111111111111111111001011000001011001110100001111111110111010,
    240'b101110011111111110111111010100101010100011111001111100011110111001111101010100010101010101010101010101010101010101010010010100100110001110000011101010011100010111010110110111101110000011001011100011100101010101010110110100011111111110111010,
    240'b101110011111111110111101011001101110100110100011011001101101001011000110010101000101010001010101010101010101010101010101010101010101001101010001010100000101001101011100011000000110000101010111010100010101001101010111110100011111111110111010,
    240'b101110011111111110111110010111101000010001011011010010001011000011010101010101110101010001010101010101010101010101010101010101010101010101010101010101010101010001010100010100110101001101010100010101010101010001010111110100011111111110111010,
    240'b101110011111111110111111010100100100111001101101101000001110101110101011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111110111111010100110100111010010000111110111110111001101011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111110111111010100010110111110000101100011101111001001110011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100011111111110111010,
    240'b101110011111111111000001010011101001001011101111110100011110101101101010010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110101001111111110111001,
    240'b101101111111111111011110010111000101100010101110110101001000110001010010010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101000001100111111010111111111110101010,
    240'b101100011111100011111110101100010110000101011000010111010101100001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100110011110111111111111111111000110101010,
    240'b110011011101000011111111111111111110010111011001110110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110011110100011111111111111111100011011010011,
    240'b111100111100100111010101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110011001100010011110001,
    240'b111110001111011011000101101011101011101111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100110110000110011001111011011110110,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule