module Background(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 600;
localparam Y_WIDTH = 430;
parameter [0:85][959:0] r_picture = {
	960'b110001101101011111011100110111001101100011000101101000000111101101011101011101101100111011100000110111111110000011100001111000101110001111100011111001001110010111100101111001101110011011100110111001101110011111100111111010001110100011101000111010001110100011100011110101111101001111011111111010001110101011101100111011101110101011100011111000011110000111011111111000101110001111100101111001011110010011100110111010001110101111101011111010111110100111101001111010101110111111110000111100001111000011110000111100001111000011110000111011111110111111101111111011111110111111110000111100001111000011110000111011111110111111101110111011011110110111101100111011001110110011101100111011001110101111101011111010101110101011101001111010011110100111101001111001111110011011100101111001011110001111100010111000011110000011011111110111111101111011011110110111001101110011011010110110011101011111010111110101111101011011010100110100111101001111010011110100101101001011010010,
	960'b011011001001011111011000111000101101111111010001101101111001010001101101011101111100100011100010111000101110001111100100111001001110001111100011111001001110010111100101111001101110011011100111111001101110011111100111111010001110100011101000111010001110010111010110110011011100111011010001110110101110010111101010111010101110100111100110111001101110010111100000111000101110011011101001111010011110101011101011111011011110111011101111111011111110111011101111111100001111000111110001111100011111000111110001111100011111000111110001111100001110111111101110111011101110111111101111111011111110111111101111111011111110111011101110111011011110110011101011111010111110101111101011111010111110101111101010111010011110100111101001111010011110100011101000111001111110011011100101111001001110001011100000111000001101111111011111110111101101111011100000110111111101111111011110110111001101101111011011110110101101101011011001110110001101100011010111110101101101001011010010,
	960'b011010000110100011101110111111001111101111111010111110001111010111110001111100011111100111111011111110111111101111111100111110111110010111100011111001001110010011100101111001011110011011100111111001111110100011101000111010001110100011101000111001111101111111010110110100011100111111010001110110001110001111101001111010101110110111101100111010111110101111101001111001011110010111100110111001101110110011101110111011111111000011111101111111011111110011111100111111011111110111111100111111001111110011111100111111001111110011111101111111011110111111101110111011101110111111101110111011101110111011101111111011111110111011101101111011011110110011101011111010111110101011101010111010101110101011101010111010011110100111101001111010001110011111100111111001101110010111100100111000101110000011011111110111101101111111011110110111101110000111111001111110111111101111111011111110111111101111111011111110101111101011111010111110101111101011111011111110001101011011010001,
	960'b100010111000011011110011111101101111010111110111111101111111100011111001111110011111011111110110111101011111010111110101111111011110011011100011111000111110010111100110111001101110011111100111111001111110100011101000111010001110100011100111111001101110010111100010110111111101111011100001111000111110101011101101111011011110110111101101111011101110111011101111111010101110100111101001111010001110101011101110111011111111000011111101111101001111010011110101111101011111010111110101111101011111010111110101111101011111010011110100111111011111000011101110111011111110111111101110111011101110111011101111111011111110111011101101111011011110110011101100111010101110101011101010111010101110101011101010111010011110100111101000111001111110011011100110111001011110010011100011111000011101111111011101110110111101101011011101110111011110000011111011111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110110111110111101011111010001,
	960'b100111101000111111110011111101101111110011110001111100011111001011110000111011101111000011110110111110111111110111110100111111001110010011100100111001001110001111100100111001111110100011101000111010001110100011101001111010011110100111101001111010011110100111101001111010011110101011101011111010111110110011101100111011011110110111101101111011101110111011101110111011111110111111101111111011101110110111101111111011111111000111111101111101001111110111111100111111001111110011111100111111011111110111111101111111011111110111110100111111001111000011101111111011111110111111101110111011101110111111101110111011101110110111101101111011011110110011101011111010111110101111101010111010101110101011101010111010101110100111101001111001111110011011100110111001011110010011100010111000001101111111011011110100101100111111011000110111001110000011111011111101011111110111111011111110111111101011111001111110101111101011111010111110101111110011110101111110101101011011010000,
	960'b101101001010001011110101111110001111000101110011011010010111000101011101010100000110000110010111110010111111101011110110111101111011111111001010110001111011110010111010110000001100101111011101111010011110101011101011111010111110101111101011111010111110101011101011111010111110101111101011111011001110110011101100111011011110111011101110111011101110111011101110111011111110111111101111111011101110111011101110111011111111000111111101111101011111110011110001111011111110111111101110111100001111000111110001111100101111110011110101111111001111000011101111111011111110111111101110111011101110111011101110111011101110110111101101111011011110110011101100111010111110101111101011111010101110101011101010111010011110100111101000111001111110011011100110111001001110010011100010110111111101111111011011110100001100110011010011110110111110000111111011111101011111101111011111110110101101001111000111110011101101011011001111110011111111100111110101111110101101010111001110,
	960'b101111111011011011110111111101111111000001011011010010010100110001000001001101110100010101011111100000001111001111111000111101001000110001101010011000000111000101111001100000011001001110100100110100001110100111101010111010101110101011101010111010101110101011101011111010111110101111101011111011001110110011101101111011011110111011101110111011101110111011101110111011111110111111101111111011111110111111101110111011111111000111111101111101011111110011101111111010111110101011101000111001111110110011101111111100011111110011110101111111001111000011101111111011111110111111101110111011101110111011101111111011101110110111101101111011011110110111101101111011001110110011101011111010111110101011101001111010011110101011101010111010001110011111100111111001101110010011100011111000101110000011011110110111001101101111011010110111001101111111111011111101011111101011010111110011101100010010111101110000001100011111000000110000111111100011110110111110101100110010111111,
	960'b011000001001000111110101111110001110110101000111010000100011100100101101001011000011011100111010010100001110111011111001111011110101010101000000010100110111001010000111100011111011011110110101100111111101001111101001111010011110100111101010111010101110101011101010111010111110101111101100111011001110110011101100111011011110110111101110111011101110111011101110111011111110111111101111111011111110111111101111111011111111000111111101111101011111110011101111111010111110100111101000111001101110011111101100111100001111110011110101111111011111000111101111111011111110111111101111111011111110111111101111111011101110111011101110111011101110111011101101111011011110110011101100111010111110101111101010111010101110101011101010111010001110011111100111111001101110010111100011111000111110001111100010111000011101111111011100110101111101010011111010111101101111100111001001110000011011111110111110101111001011101010111000110000001111100011110110111110001100000010110111,
	960'b001001110011111111101101111110101110101100110110001011110011010100100001001001000011001100110011010001101110110111111001111011100101100001011110011011101000111110101011101100011100010111011101110010101100001111100100111010011110100111101010111010101110101011101010111010111110101111101100111011001110110011101100111011011110110111101110111011101110111011101110111011101110111111101111111011111110111111101111111011111111000111111101111101011111110011101110111011001110101011101001111001111110011111101100111011111111110011110101111111011111000111110000111100001110111111110000111100001110111111101111111011101110111011101110111011101110111011101110111011011110110011101100111011001110101111101010111010011110011111100010111000111110011011100110111001011110010011100100111000111110001011100001111000011101111111011000110011011100101011111001111101101111100111000101101111111100000111000001101110111011100110111001101110101111100011110110111110001100001111000000,
	960'b001000000011000111101011111110101110110000110101000110010010000000011110001000010010100100101001001111001110110011111001111011100101110101110010100011011010101111001010110110101101110111100101111010001110001011100110111010011110100111101001111010101110101011101011111010111110101111101100111011001110110011101101111011011110110111101101111011101110111011101110111011101110111111101111111011111110111111101111111011111111000111111101111101011111110011101110111011011110110011101010111010011110100011101100111100001111110011110101111111011111000111110000111100001111000011110000111100001110111111101111111011111111000011101111111011111110111111101011110111111101110111100111111001101110100011101001111001101101011111001000110010111101110011100100110110111101001111011011111000011110001111100000110111011101100011001011101111111100010011111001111101101111100111000101101111111011111111000000101110011011100010100110100101011111001111110111111110011100010111000011,
	960'b010011010100100111101101111110101110101100101011000101000001100100011110001000000010010000100100001111011110110111111001111011110110010101111100101011001100110011011101111001011110011011100111111010011110100111101001111010011110100111101010111010111110101011101010111010111110101111101011111011001110110011101100111011011110110111101101111011101110111011101110111011101110111111101111111011111111000011110000111100001111000111111101111101011111110011101111111011111110111011101100111010111110101111101110111100001111110011110101111111011111000111110000111100001111000111110000111100001111000011110000111011111110101011100110111010101110110111011101110011001101001111010101110011011101100011100010110111011100100110111101101111101100110111011000110010101100010111000111110100001110000011011101110100001100100111000010101111001100001011111000111101101111100111000101101111111100001111000100101110101001001101100010011110101111001011110111111110011100101111000000,
	960'b100011110111110011110001111110011110101100101000000100010001100000011101001000100010001100100011001111011110110111111001111100100111101010001101110001101110000011100111111001101110011011100111111010001110100011101000111010001110100011101001111010101110101011101010111010101110101111101011111010111110110011101101111011011110110111101110111011101110111011101111111011111110111111101111111100001111000011110000111100001111000111111100111101011111110011110000111011111110111111101110111011101110111011101111111100011111110111110101111111011111001011110001111100011111000111110000111100011111000111110001111010001101010111010000111000001110010011010101110010101100100111000101110001011100100111001001110001111100000010111100101111011100010011001001110001101100001011000011110011011101100011010100110001111100000011000000101111101100001111111000111101101111100010111111101111011100001010111111101010100101100101001011011110001111001111110111111110011100011110111100,
	960'b011011010111011111110001111110011110111001000100001011000010111000111011001110100011010100110110010010011110111011111001111011110110010101110111101100011101010011100011111010001110011111100111111010001110100011101000111010001110100111101010111010111110101011101010111010111110101111101100111011011110110111101101111011011110110111101110111011101110111111101111111011111110111111101111111011111110111111110000111100001111000111111100111101011111110111110010111100011111000011110000111100001111000011110001111100101111110111110101111111011111001011110001111100011111000111110001111011101110111111110000110111101100111111001100110100111101010011001101110010001100001111000000110000011100000110111111101111111011111111000010110000111100001111000010110000101100011011001100110011001100101011001010110000101011110110111101101111101100001111111000111101101111011010101011101110011100000110111100100101100101011101011001100001001111010011110111111101111011000110110000,
	960'b000111110011010111101100111101111111101111101101111010111110101111101101111011001110110011101100111011011111101111110111111011100101100001010100011010010111110010100010110011101101111111100111111010011110100011101001111010011110101011101011111011001110101111101001111001101110001111101001111011001110110111101101111011011110110111101101111011101110111011101110111011111110111111101111111011111110111111110000111100001111000111111101111101001111110111111101111111011111110011111100111111001111110011111101111111011111110111110100111111011111001011110001111100011111000111101100110111011110011011101101110111001101001011010000110011001100100111001010110011001100101111000101110001011100010010111111110000011100001111000110110001011100000010111111110000101101000011010011110010111100100111001001110000011011111010111111101111111100011111111001111101011111110011110110111101111111100011111000111101001110111111101111111100111111110011110101111101101010011110101010,
	960'b001000110011100011101110111110011111011111111001111110101111101011111010111110101111101011111010111110011111011111111000111100100110010001100111011111110111101101111001100110001011110111010001111000111110101011101001111010011110100111101010111010101110101011100011110110101101100011100011111011001110111011101110111011101110111011101110111011111110111111101111111100001111000011110000111100001111000011110000111100011111000111111101111101001111010011110101111101011111010111110101111101011111010111110101111101011111010011110100111111011111001011110001111100011110110011100010110100111101111011101010111000101101101011010010110011011100100111001011110101111101111011001110110011101100110111000001110000101100001011000011110001011100000111000000110001111101010011010000110001111100010111000110110001001100000111000001110000101100101111111100111101111111011011110111111101111111011111110111111110001111100111111001111110001111011111110111111101111010010110100011,
	960'b011000100111011011101010111011111110110111101111111011101110110011101011111010111110101111101101111011011110110111110000111001110111100101101011011011010110111001110110100010111010101011001001110011001110000111101011111010011110011011100011111001101110100111100000110101101101010011011011111010001110101011101101111011101110111011101111111011111110111111110000111100001111000111110000111100011111000111110001111100011111001011111101111111011111110111111101111111001111110111111101111111011111110111111101111111011111110111111101111111011111001111110000111010011101110111010100110101111110010011101101111011001110001111011100110101011100111111010010110110111101011111001100110001111100011111000010110000101100000111000010110001001100000010111110110000111100101111000101110000001100000111000010101111111011000110011101100011111001010111100111111100011111010011110100111100011110111111110000111011101110110111101111111011111111000011110010111011111010011010011001,
	960'b101001111001110001111100010010000100000001001111010001100011010000101011001010110010111101000001010001110100100001011000011001000111100010010101100100100111111001110000011011011000101011001100111000001110000011101000111010011110000111011011110111011110000011010110110101011101011011001101110011001101110011100011111010111110111111101111111011111110111111101111111011111111000011110001111100011111000111110001111100011111000111110010111100101111001011110011111100101111001011110010111100101111001011110001111100101111001111110011111100111111000111101001110111011101011111010111111000101110111011110001111100101110110111100111111000011101101111010111110100011100100011000100110000101100001011000011110000101100000111000010110000011011111110111110110000001100001010111110101111101011110110111110101100011000110001101101010101000100011101001110010111111000000010000101011011000101011001011110010010110100010001010001010110100101111001110010100101101001100110100010,
	960'b010110100011110000100100001000000001111100100100000111010001100100011010000110010010001100111101010011010100001101001001010011100100011001011011100001001001110110100101100110100111101110101000111001011110100111101001111010011110011111100010110110111100110110111001101110111101000010101001101000111100011111000001110111101111000011101111111011111110111111101111111011111111000011110001111100011111000111110010111100101111001011110010111100011111000111110001111100101111000111110001111100011111000111110001111100011111000111101111111011111110101011100010110111011101110111011111111001011110111011110000111100001111000011101100111010001101110011001001110000111100011011000100110001011100001110111110110000001100010111000100110000101100000010111111110000001100000110111110101111101011110110111100101101011010101110100100100110010111111001010111001101000010110101000011010101000100001000111000001011110010111000111001001111010100100101101011100000101001010010011100,
	960'b000111100010000100101000001100110011001100101011001000100010001000100010001000010011001101001000011000111000000101111100011111010110001001010011011000010111111010011100101110111010100001111111101110111110010011101000111010001110011111100100110101011011100110100011100110011011001110011001100011111010001010111110111001011111000011110000111011111110111111110000111011111110110111110001111100011111000111110001111100101111001111110011111100111110110111100101111010111111001011110010111100011111000111110001111100011110111111101101111011101110110111100111111001101110100011100101111001101110100111101000111010001110101011101011111010001101101010110111100000011001001110110110110000101010101110010001101010001100100111001000110001011100001111000011110000101100000010111111101111101011111010111101101111011011110010111111101100111000101101101010010011100010111000011110001001100010110100100111001001010010110100111000001110010100110001101001011110010111111101110101,
	960'b001010010011010001000001010100010011100100100011001001010010000000011110000111110100001001101110010100010110011101111100100001101001001101111001010111110110011110001100101100111100011110100100100110001100011011011101111000011110001111011100110100011100011010101101100010110111111001111000011100001000010010100001101111011110000111110000111011001110101111101000110111011101100111101001111011011110000011100000111011011111001111110011111010111101001011000000110001111101110111110000111100011111000111110001111100011111000111110001111100011111000111101111111011111111000011101101111010001110011111100100111000001101111111100100111001101101111010110111011100000100111101100111100011100110101001101000101010001100100110110110101110101100010111000011101111011011110110111111101111111011111110111111101111101011110110111101101011011010001010010001011101000100011100101001000110110001100000011001000111100010011100101110001100100100110001101011011001000100010000111000,
	960'b010011000101101101100000010111100010111000100001001001100010001000100001000111100100011110010011011011000100011101110101011111001000111110011110011111010101101101110001101011011101000011010110110001111100001011001011110101001101010111010011110011101100010010101100100011110110110101011110010111110111000110010001101011001101000111101011111010101110011011010110110011101100101111010101110110111101011011011110111011001111001111110010110110111011100110110000101100101011111111011111111011111111000111110001111011101110111011110001111100101111000111110000111100001110111111101111111011011110110011100100110000011010101010111011110110001110000011001010100011100100101000111011010100110100111001100001100110011001110001111111101011011011110110101000100111111010111110111101110000011100000010111111101111011011110110111101101111011100001010111100101001000111111101010101001010100001100100010110000101110001110000100010001010110011100100110101001001100010010000101110,
	960'b011100000111110101110000010010100010001100100110001010100010101000101010001001110101011110011011011110010011111001001011011111011000010010010011101010000111101101011011100101111101100111100001110110111101011011001011110100001100101111001001110010011100000110101101100011010110011101010110010110000110100010010011110100101110010011101000111001111101111111001001110001101100011011000111110100001110000111101110111011111110011011100100110010011010111010101110101110001011110011000011110111011110100111011000110011001100111111011111111100011111000111110000111011111110111011101101111011011110110011101001110110011011001110001110100100101011110011001000100100110100111000110100001110100011111101001110011010110110110101111011100101101000010010000010100111001011101011000010110000011100000010111111101111011011110110111010101110101011110110111101101101111001100101101100010000100010010000011000000101100001100000101001001101000010001000011101001001100011000000111100,
	960'b100010101000010101010111001001010001111100101110001101100010110000101100001111101000011010100001100000000101001100110111010100011000110010010010101011011011001001110111011111111101010111100011110110011101000111010001110101011100111011001000110010011100100110111010100100100111100101010110010011010110101101111110101100111101001111011101111000111101000111000001110000001100000111000110110100111110001111101000110110011011111010111001101100111010101110111000110010101011110010110000101111101100011010110100101100001011011011010000111011111111001011110000111100001110111111101111111011111110110111101011111010011101101110110110100100101000001110011011100110110101000100101110001100110100000001000010010011100110011101101011010100110101111010001111101111011101000011000110110000101100000110111111101111111011110010111001101110001011100110110100101001101001010001111010010110100011000100100000000110110001111001000100001101000001111000101100010010010101010001010100,
	960'b100011000110101100101110000111000010010000110111010001110010110000101010010110111001100110011110100011010111001101010000001101000101110110011011101001001100100010110010100010011011111111011010110100001100101011001010110011001100111011001011110011001101000011000100100110100111011001010110010010100110011110010001101000111011100110111111110000101011101010110111101101101011100010111101110011001101001011000001101011111010101110101011101011001010110110110110101110111011001010101111101100011011001010110000101100011011010011000111111001011110110111101011111001001110001011100001111000001101111111011101110111011101110011000110101100001001101001111001011101110101110000111001001110110011111101000001010011000101011101000000010001100110101010011000101111011100101011000101110000111100001011000000110000001011110110111011101110111011101010110001100110001000001001110001010111110100011100110000001001010010010000110011001000110010011100110111001111110100011001001010,
	960'b011001010011100000011110001000110011001000111111010011110010111100101111011100011001000110010001100011011000100101101011001110100011100101101100101000101100001011010000101100101010110011001001110010001100011111000110110010001100110011001000110010011100101010110001100010011000001110000011100000000111111010000001011111100111101001110111011100100111000001101111011011010110111001101011011011000110101101100111011100111010000110111011110001011100110111010110111000111110100011101100111011011110110111101010111000111101011011001110110010011011111110101010011110110110101101101010011010000110100101101010011100010111011001111000011110000111101101110110011110010111101001110101011100100111001101110000011100010111000101000001010101110111011110011111110000111100101111001011110010001100001111000100110010001100000110111100101110101011011110101011100010010110010001001110010000010011000000011110000101110001100000011000000110100010011000101110001110010100010101001011,
	960'b001110100010001100100001001100010100011101010001010100010010110000110111011111001000110010001100100011101000101101111100010100010011010101000101100001011011001011001000110010001011001111000000110000101100000111000010110000111011110010010000100010101000110110010011100100101001000010001101100011011000100110000100011111000111010101101111011010000110010001100011011000110110001001100001011000110110001101100000011000000110100110010100100111101010001010100100101010101010110010101111101011111010111010101101101010111010010110100001100111001001000101101000010111000110000101100010010111110110000001100000011001110110110001101110011100000111001101110111011110100111110101111101011111010111111010000000011111100111100101101111011111000111100110000001100101111011001011000110110010011100011111001110110100001100011010111011101101101001011001100000010000110011011000110000001011100010011000010111000101010001011000010011000101010001011000011101001101100101010001011110,
	960'b001001010010001000101111010001010101100101100101010110000011000101010100100000111000100110001010100011111000110110000100011001110011111101000010011000001010001010111011110000111011001010111000101111101011110110110111101100101000011010000101100100001001100010011111100111111001111110011010100101111001000010001100100010001000100110000110100000010111111101111111011111000111100001111000011110000111100101111000011110100111100101110111011101100111011101110101011101000111010001110100011101000111010001110101011101100111011101110110011101100111010101111011011110010111101001111101011110100111101101111000011110100111111001111111100000111000011010001001100010101000101110001010100010111000100110001101100100001000111010000101011111000111010001110001010100100111001010100111110010001101000111010100110100011100011110111000100101000101000100110110001111010101000101011011010000010011001000011111000111010001110000011011001001100001111000010111000111000011111001101000,
	960'b001001110010110100111111010100100110011001110001011001110100010001110100100001001000010110001001100010111000101110001000011111010101001001000110010100011000001010101111101110011011001110110111101110001010110110000000100001001001010010100101101110111101001011100101111001101110001011011011110110011101100011011000110101101101011011010110110101011101010111010101110101101101010011010101110101101101011011010111110110001101100011010110110101011101010111010101110101011101010111010101110101001101010111010101110101011101010111010101110101011101010111010110110101101101010111010110110101011101010111010100110100101101001111010011110100111101001111010100110101011101010111010101110101011101100011100000111001011101111111000001101001001000111110000011011101010111000101111010101111001101011011010001110011011100010010011010010101010011100001000110011010111000100101110111010000010010111000011100000110000001100000100101010001000011010000100110000110010001101000101010,
	960'b001100010011111101001100011000010110111001110101011011000101001110000000100001111000010110001001100010111000110010001011100010010110100001001100010100010110110110011011101010011010111110110010101010001000101110001010100110001011101011010101111000001101100110110111101001001001101010010010100100011001001010010010100100101001000010010001100100101001001010010010100100111001001010010010100100101001001010010010100100101001001010010001100100101001001010010010100100111001001110010011100100101001001010010011100100111001001110010011100100111001001010010010100100101001001010010010100100101001001110010011100100011001001010010010100100011001000110010001100100011001001010010010100100101001010110100001101100101100011111100010110111011100010110100111100100011000100010001000101011011100100011001101110011101011000001011100001111000100101001101110100101001001100001111101010010110010101000011001000101110001100100101101010111000101101001000101001100110001111100011001,
	960'b001110010100111101011100011011000111010101110100011001000101100110000101100100001000111010001011100011101001001010010001100011000111101101011111010110010111000110001010100110101010000110100100101010001010010111000100110110011011010110010011011101100101000100011110000100010000111100001110000011010000110100001101000010110000101100001011000010110000101100001011000011000000110000001100000010110000101100001100000010110000110000001100000010110000110000001100000010110000101100001100000011100000110000001100000011010000110000001100000010110000110000001100000010110000101100001011000011000000101100001011000010110000101100001100000010110000110000001100000011000000110000001100000011100000110100010001000110010010111101101111100100001011000011010011110100101011010110110011101100011011101111000111101111000110111101000010010101010111011110011001101000101001101010001110010101110011001100011101000110110010000100110010011001000111100001101101010111100011100100100011,
	960'b010001000110000101101100011100100111011001110010010100100101100110001001100110011001110010010000100011101001000010010000100011001000100101110101010111000111101110001110100101101010100110110101101011101100110111100001110001100111000000111010000101100000011100000011000000010000000100000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000010000000100000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000010000000100000000000000100000001000000010000000100000001100010001001100110110010110010111111000011101111111000011101111111011011110111010100011110101001001011001100000001001111010110101101101011011000110011000010100110010100100011110000111100010011100110110011000101000001110000010011101000101101000111111,
	960'b010101010110110001110011011100010111001101101100010000110110010110001110100101111001010110001010100000111000010110000110100001001000010101111101011000110111011010010010101001111011011011000000110010101101010010110001011110100001101100000100000001000000001100000100000000100000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000001000000010000000011000000110000001100000011000000110000010000000100000001000000010000000011000000110000010000000011000001000000010000000011000000110000001100000011000000100000001100000100000000110000010000000011000000110000001100000011000000110000001100000100000000110000001100000011000000110000010000000011000001000000001100000011000000100000001000000011000001000001000000111110101000111101100111011100110001011100011110110110100111110110011110001001101001001011010110111110110000001011110110010111010000100010001100100101001000100010111001000110011011111000100110001001011111010110111001011000,
	960'b011000010110110101110001011011110111000001100001001111010111010010000100011111110111110001111100011111000111111010000000100000011000000110000000011101000111101110010001101110001011000011000000101010100110010100100000000010110000001100000010000001000000011000000010000000100000001000000001000000100000001000000001000000010000000100000001000000100000000100000001000000100000001000000010000000100000001000000001000000010000000100000001000000100000001000000010000000010000000100000001000000100000001000000001000000010000001000000010000000100000001000000001000000010000001000000010000000100000001000000010000000010000000100000010000000010000000100000001000000010000001000000001000000010000000100000010000000100000001100000101000000110000001000001000000110100101100010100010110101111011111011000110101110001000110110101001101100001011100110111011101111111011110110001101001101010010101000110110001010000011011001010101011110101000100010001000011111110111001101101000,
	960'b011001110110110001101110011011100110110101010001010000110111000101110110011101010111100001111001011110010111110001111101011111100111111110000000011111100111111010010001101010111011101011000110011000000001010000000001000000010000001100000110000001100000001000000001000000010000000100000010000000100000001000000010000000100000001000000010000000100000000100000001000000010000001000000010000000100000001100000001000000010000000000000001000000010000000100000010000000010000000100000010000000100000001000000010000000100000000100000010000000010000000100000001000000010000000100000010000000100000001000000001000000010000000000000001000000010000000100000001000000100000001000000010000000010000000100000010000000100000000100000100000001010000010000000011000000100001000001001101101000001100111110111100101111011000110001111010101010101011001110110101101100111010111001110011001100000011100101001001001011100100001101100010011111111000010010000100100000100111101001110010,
	960'b011010100110101001101011011011010110100101000010010100000110111101110001011100110111010101110111011110010111100101111011011111000111110101111110011111010111100010001100101111011100100001111010000100000000000000000010000001000000001000000011000000100000000100000010000000010000001000000010000000100000000100000001000000100000000100000001000000010000000100000010000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000001100000010000000010000000100000010000000100000001000000010000000010000001000000001000000010000001000000001000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000100000000100000001000000100000001000000010000000100000001000000100000000110000001000001000001001101100001111011111101101111000010101111000101000101010101110101001101000001001000001010100001101100101010001101000001101100100110001110000100000011000001010000010100000100111110101110100,
	960'b011010010110100101101010011010110110001000111101010111110110111101110001011100110111010001110100011101100111100001111011011111010111110101111100011001100111001110001100110000111001011100110001000001000000001000000100000001100000001000000001000000100000000100000001000000100000001000000001000000100000000100000010000000010000000100000010000000010000000100000001000000010000000100000001000000010000000000000001000000010000000100000001000000010000000100000001000000100000001000000001000000010000000100000010000000010000001100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000000000000010000000100000001000000010000000100000001000000010000000100000000000000010000000100000001000001010000001100000000000011001000010111011000110011011000001001101111011100111001110110010111100100001000000101000110010000100110101001110111010000110101001101111010100000001000000010000001100000011000000001111100,
	960'b011010010110100101101010011010100101010001001000011011000111000101110010011100110111001101110100011101010111100001111010011110110111110001110111011000010111011010011110100010110010001100000101000000100000010100000011000000100000000100000010000000110000001000000010000000010000000100000010000000010000000100000001000000100000001000000011000000100000001000000010000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000001000000010000000010000001000000010000000100000001000000001000000100000000100000001000000010000001000000001000000100000001000000010000000010000000000000001000000010000000100000001000000010000001000000010000000010000000100000010000000100000001000000010000000110000001000000010000000100000010100000011000000110001101001111011110011111000101001100100011001011001000110010000100010100110110100111100010100000111010101111011010011010101110010000000100000011000000010000001100000011000100110010101,
	960'b011010100110100101101010011001110100010101001101011011110111000101110010011100100111001001110100011101010111011101111001011110110111100101011011010111101000001110101000010011000000011100000010000000110000010100000001000000010000001000000010000000100000001000000001000000010000001000000001000000010000001000000010000000100000000100000001000000010000001000000010000000010000001100000010000000010000000100000001000000010000000000000001000000010000000100000010000000010000001000000001000000010000001000000001000000010000001000000010000000010000001000000001000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000010000001000000010000000010000000100000001000000100000000100000010000000010000001100000011000000010000001000000110000001000000010000110111101100111001111001100101010110100110000010000111100010010110000001000010011000010111101101111100010100010101101101111111100000011000000110000010100001101000111010010101,
	960'b011010100110100001100110011000010100010101100000011011110111000001110001011100100111001001110101011101100111011001111000011110110111100101010111011001011001010110101110001000110000001100000011000001010000001000000010000000010000001000000001000000010000001000000001000000100000001000000001000000010000001000000010000000100000000100000001000000010000001000000001000000010000001000000001000000110000000100000000000000000000000000000001000000010000000000000010000000010000000100000000000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000000100000001000000010000001000000010000000100000001100000010000000010000000100000001000000010000000100000001000000100000000100000001000000100000001100000010000000100000000100000101000000110000001100010100011111011010111101110011010101110101100110000101100001000101101001010001011011100111110101111101010100010101001001111111100000101000000110000010100001111000101010001011,
	960'b011010010110010101100100010110010100010001101000011011110111000001110001011100100111001001110100011101000111010001111000011110100111010001011001011101111010101110101000000100100000000100000100000000110000001100000001000000010000000100000010000000100000000100000001000000010000001000000001000000100000000100000001000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000000100000000000000010000000100000010000000010000000100000001000000010000000100000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000000100000001000000100000001100000010000000010000001000000010000000100000001000000010000000010000000100000001000000010000001000000001000000010000001000000011000000100000001000000010000001100000010000000100001010101011011010010001010111000101011010000100100000110110011001100101011110000111111101111110010110000100101001111110100000011000000010000010100001011000101010001111,
	960'b011010010110011101100100010011000100011001101100011100000111000001110000011100000111000101110011011100100111001101111000011101000100101001011001100001011011001010001111000011100000000000000100000000100000000100000010000000100000001000000010000000100000001000000001000000010000000100000001000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000000000000001000000010000000100000001000000010000000100000001000000100000001000000001000000010000000100000001000000010000000100000010000000100000001000000001000000010000001000000010000000100000000100000001000000010000000100000001000000100000001000000001000000010000000100000010000000100000001000000010000001010000001100000010000101011011011110011111011001000101011110000001100000100111010001111000011111010111111101111111011000000100001101111101100000101000000010000001100001001000110010010001,
	960'b011010000110100101100100010000010101001101110010011100110111001001110010011100100111001101110100011100100111011001111001011101000100100001100101100101111011001001011001000010010000001000000101000000010000001000000010000000100000001000000001000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000000100000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000001000000001000000010000001000000001000000010000001000000001000000010000000100000010000000010000000100000010000000010000000100000010000000100000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000110000001000000010000000110000010000000001000100011010111010101001011101010101110001111111100000010111101101111110011111110111111101111111011001100011110101111000100000100111111110000000100000011000010110000101,
	960'b011010010110100101011111001110010110011101111010011110010111011001111000011110110111100101110111011101010111100001111010011101000100110101101101100111011010111001000001000001110000000100000100000000100000000100000001000000100000001000000010000000010000000100000001000000010000000100000001000000010000000100000001000000100000001000000010000000100000001000000001000000010000000000000001000000100000001000000001000000010000000100000010000000100000001000000001000000010000000100000010000000010000001000000001000000010000000100000001000000010000001000000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000000100000001000000010000000100000001000000010000001000000010000000100000001000000010000000010000001000000001000000100000001000000001000000010000001100000010000100001010010010101010011110110110000101111111100000100111111101111111011111110111111110000000011011000011100101110011100000010111111101111111100000001000000110000001,
	960'b011011000110110101010111001111100111111010001010100001010111111110000000100001101000010001111101011110110111110101111100011101000100111101110010100111111010100100110101000001010000001000000101000000100000000100000010000000100000001000000001000000100000000100000010000000010000000100000001000000010000000100000001000000100000001000000010000000100000001000000001000000010000000100000001000000100000000100000010000000010000001000000010000000100000000000000000000000010000000100000001000000010000000100000010000000010000000100000010000000010000000100000001000000010000000100000001000000100000000100000001000000100000000100000010000000010000000100000010000000010000000100000001000000010000000100000010000000010000000100000001000000100000001000000010000000100000001000000011000000100000001100000010000100011001101010101011100000100110011001111111100000011000000010000000011111110111111010000000011100010011011001101100100000011000000101111111011111110111111101111110,
	960'b011101100111011001001011010011001000010010001001100001101000010110000011100001001000010010000001100000000111111001101111011000100101001001111010101000001010010000110000000001000000001000000101000000100000001100000011000000110000001000000010000000010000000100000001000000100000000100000001000000010000000100000001000000100000001000000001000000100000001000000011000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000100000000100000010000000010000000000000001000000010000001000000000000000010000000100000001000000100000001000000010000000100000001000000010000000010000001000000001000000000000000100000010000000100000000100000001000000100000000100000010000000010000000100000001000000100000001100000001000100011001000110100110100001100110111110000000100000101000000110000000011111110111111110000001011101010011100001100100100000001000000001111111011111100111111001111101,
	960'b100001110111101100111101010110111000000110000010100000011000010010000100100001001000001101111111100000000111001101101010011010110101100001111111100111101010010100111000000001100000000100000100000000100000000100000011000000010000001100000010000000100000001000000001000000100000000100000001000000010000000100000001000000100000000100000001000000010000000100000010000000010000000100000010000000000000000100000001000000010000000000000001000000010000001000000001000000010000000100000001000000010000000000000000000000100000000100000001000000000000000100000001000000010000000100000000000000010000000100000001000000010000001000000010000000110000000100000001000000010000000100000001000000010000000100000001000000100000001000000010000000100000000100000010000000110000001000000010000000100000010000000010000100011001010110100010100010010111011010000001100000101000001010000001100000000111111110000001011110010011110001011001011111110111111101111110011111010111111001111101,
	960'b011111110110101100110111011011011000001010000010100000001000001110000110100001001000001101111111100000100111101010000001100000000110010010001110100110011010101101010101000010110000001000000101000000110000001000000010000000110000001000000010000000010000001000000010000000010000001000000001000000010000000100000000000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000010000000010000000100000001000000010000000100000010000000010000000100000001000000000000001000000010000000100000000100000001000000110000000100000001000000010000001000000001000000010000000100000001000000010000000100000010000000100000000100000010000000100000001000000010000000100000001000000011000000110000001000000010000100101001110110011100100110001000010010000011100000111000001010000010100000010111111110000001011111000100000101001101011111101000000001111110011111010111110101111101,
	960'b011101000101001100111011011110101000010010000100100000011000001010001000100010001000010110000011100010101000100110001010100001110110101110011001100110101010101101101110000011010000000100000100000000110000001000000001000000010000001000000011000000100000001000000001000000100000000000000001000000010000000100000001000000100000000100000001000000010000001000000001000000010000001000000001000000010000001000000001000000010000000100000001000000010000000100000010000000010000001000000011000000100000000100000010000000100000000100000010000000100000001000000001000000010000000100000010000000010000000100000001000000010000000100000001000000010000000100000010000000010000001000000001000000010000000100000010000000010000000100000010000000100000001100000010000000100000001000000011000001000000001100000011000100101001111010011011101001101001000010000111100001001000010010000011100000101000001010000001011111100100110001000010011110100111111101111110011111010111110101111101,
	960'b011011100011110101001100100001101000101010001010100010001000010010001011100011011000011110001000100100001001000110010010100011100111001010100110101001001010011010001000000100010000000100000010000000110000001000000001000000010000001000000010000000100000001000000010000000010000000100000001000000010000000100000001000000010000000100000001000000010000001000000001000000010000001000000010000000010000001000000001000000010000000100000010000000010000001000000010000000100000001000000010000000100000001000000001000000010000001000000001000000010000001000000010000000010000000100000001000000010000000100000001000000100000000100000001000000010000001000000010000000010000000100000001000000010000000100000010000000010000000100000010000000010000001000000010000000100000001000000011000001010000010000000100000110011001110010011111101101101001110110001100100010101000011110000111100001011000010010000101100001000101100100110111011101100111111101111110011111010111111001111101,
	960'b011000100011001101101000100011111000111110001110100011011000011010001110100011111000100010001111100101111001100010011001100001100110100110110110110001101001110110011101000101000000010100000100000001010000001100000001000000010000001100000010000000100000001000000001000000010000000100000010000000100000000100000001000000010000000100000001000000100000001000000001000000010000001000000010000000100000001000000001000000010000000100000001000000100000001000000010000000100000001000000011000000100000001000000010000000100000001000000010000000100000000100000001000000100000001000000010000000010000000100000010000000010000000100000001000000100000000100000001000000010000001000000010000000010000000100000010000000010000001000000010000000100000000100000010000000100000001000000011000001000000010000000111001111111001000110111101110001111010111110010010100011111000110110001011100010101000011110001000100001110110011100110001011100011000001001111111011111111000000001111110,
	960'b010011100011111010001101100111111001110110011100100110111001011010011100100111101001010110100001101001111010100110101011100011110101101010110101110100101010101010011000001000100000011100000100000001010000001100000001000000010000001000000010000000100000001000000001000000100000000100000001000000100000001000000010000000010000000100000001000000010000000100000010000000100000000100000001000000010000000100000001000000000000000100000001000000100000000100000001000000010000000100000001000000100000000100000001000000010000000000000001000000010000000000000001000000100000001000000010000000010000000100000010000000010000000100000001000000010000000100000001000000100000000100000001000000010000000100000010000000100000001000000010000000010000000100000010000000110000001000000101000000110000010100010110011011101001101011001111110010101011010110011000100101001001001110010010100100001000110110001011100010110111001100110001011010001000010010000011100000101000001010000010,
	960'b001100000101101011101001111101101111010111110101111101011111010111110101111101011111010011110110111101101111011011110111111010010111110110110001110010101100111010011010011100100001100000000101000000110000010000000101000000110000001000000001000000000000001000000010000000110000001000000001000000010000001000000001000000010000000100000001000000100000001000000010000000010000000100000001000000000000000100000001000000010000000100000001000000010000000100000010000000010000000100000010000000100000000100000001000000010000001000000011000000100000000100000010000000100000000100000000000000000000000100000001000000100000001000000010000000010000000100000001000000100000001000000010000000100000001000000010000000010000000100000010000000100000001100000100000000110000010100000011000001000001000001101000101001101100101011010100110000001010001010011111100111011001110010011011100110001001011010010010100011110111110100110010010111001000011010000111100001111000011010000110,
	960'b001010100111110111110110111101111111011011111000111110001111100011111000111110001111011111110111111101101111010111110110111101111010100110101110101110101100011110110101100111110100101000001010000000110000001000000100000000110000001000000001000000100000000100000010000000110000001000000010000000010000001000000010000000010000000100000001000000010000000100000001000000000000001000000010000000010000000100000000000000010000000100000010000000100000001000000010000000100000001000000010000000100000001000000001000000010000001000000011000000100000000100000001000000010000000100000000000000010000001000000010000000010000001000000010000000100000001000000010000000100000000100000010000000100000001100000010000000100000001000000010000000100000001000000010000001010000001100000100000001110011010110010111101000111101010111000111101101101000001110101000101011001010100010100111101001001010001010011110100110111000101100111010010011101000011110001010100010001000100010000111,
	960'b001100110110101111110010111101101111101111101110111011011110110111101101111011111111010111110111111110101111110011110101111110101100010110001010101001001011000010111001101001001000101000101101000001010000001100000100000001100000001100000001000000010000001000000001000000010000001000000010000000100000001000000001000000010000000100000001000000010000000100000001000000010000000100000010000000100000001100000010000000100000001000000011000000100000001000000010000000110000001000000001000000100000001000000010000000100000001000000010000000100000000100000010000000010000000100000001000000010000001100000010000000100000001100000010000000010000001000000010000000010000001000000001000000100000000100000001000000010000000100000010000000010000001000000010000001000000001100000011000100100111100010100001100101011100000010110010101001011010111010110100101100111010111010101100101010101010011110100110101000101001010101001001010001001000010110001010100010101000100110001000,
	960'b001011010011111111101101111110101110111001001110001111100100010101000101010100011000100110011010101110101111100011110110111111001100100001000100011100101000110110001101100011101001011010010001000101100000000100000011000001000000010100000101000000010000001000000010000000010000001000000001000000100000000100000001000000100000001000000010000000110000000100000010000000100000001000000010000000100000001000000011000000100000010000000011000000110000001000000010000000010000001100000011000000110000001100000011000000110000001000000011000000100000001000000011000000100000000100000010000000100000001000000010000000100000001000000010000000100000000100000001000000100000000100000010000000010000001000000001000000100000001000000010000001000000010100000100000000110000001000001001010001011001001110010100101010101001101010001010010101111010000010101010101001111010000010011010100110001001011010010100100100101000110101010111001111011000000010001010100010101000100110001000,
	960'b001001010011011011101100111110101110110100111110001011010011000100110000001100110011111100111100010110101111000011110111111110101101100010111011010001010111000101110111100000101000010010010101010100010001010100001010000001000000001100000101000001100000010100000001000000010000001000000010000000110000001000000010000000100000001000000011000000100000001100000011000000110000001000000010000000100000001000000011000000110000001100000011000001000000001100000011000000100000001000000010000000110000010000000010000000100000001100000010000001000000001000000011000000110000001000000011000000100000000100000010000000010000000100000010000001000000001000000011000000100000001100000011000000100000001000000010000000010000001000000110000001100000001100000011000010000001000100111100100011111000100110010110100101101000001001100001100010101001011110011000100101111001011010010101100100111001001010010010100100011000111101101010001101100111011010001010100010101000101010001000,
	960'b001000000011010111101100111110101110110000111001001010110011001100101111001011000010101100101001001111101110110111110111111110101101111111001111001111010010100001010100010111100110010001110101100101111001100001100011000111010000010100000100000001000000010000000011000001010000010100000100000001000000010100000100000001000000010000000100000001010000010100000100000001010000010000000100000001000000010000000100000001000000010000000101000001010000010100000100000001010000010100000100000001010000010000000101000001010000010100000100000000110000010000000100000001000000010100000101000001010000010000000100000001010000010100000110000001010000010100000101000001010000010000000100000001010000010100000101000001010000001100000100000000110000000100001001010100001001010010011010100010011000000101111011011100000011111100110110100100001001100110010111100101101001011010010110100100111001000110010001100100001001000001111010001101100110100110001001100010101000101010001001,
	960'b000111110011010011101100111110101110110000110101001001000010100000100101001000010010000000100100001110101110110011110111111110111110001011011111110001110011101100101101010011010101100101100000011110011001100110100001011101010001101100010000000011010000100000000010000001000000010000000011000000100000010000000100000000110000001100000011000000110000001100000011000000110000001100000011000000110000010100000011000001000000010000000101000000110000001000000100000000110000001100000011000000110000001100000011000000110000001100000100000000110000001100000011000000110000001100000100000001000000001100000011000001000000010000000100000001000000001100000010000000110000001100000100000000110000010000000010000000110000010100001101000100010001000000101110100111001010000110000111011111100111100001101110011000110011011110000111100110101001100110011000100101111001011010010110100101011001001110010010100100011001000110000100001110010101010110001001100010111000101010001010,
	960'b001000010011010111101100111110101110110000110111001001100010011100100000000111000001110000011100001101001110110011111000111101101010001110010100110010111100101100111111001101010101000001001111010110000110010101110100100001001001101010001110011000110011010100010000000010100000100100001000000001110000011100000111000001010000010100000100000001010000010100000111000001100000011000000111000001110000011000000110000001110000011100001001000001110000011100000111000010000000100000000111000001110000011100001000000001110000011000000110000001110000011100000101000001010000011000000110000001010000011000000110000001100000010000000101000001100000011000000111000010000000100100001000000010000000100000001001000011000001111101101100100101011010000010010110100010011000001001110100011011100110101101010010001111101000101110011101100110101001100110011001100110001001011110010111100101111001011110010100100100101001001010001011010001000100011010000110100010111000101110001010,
	960'b001000110011011111101100111110101110110000110101001000110010100100100110001000010010000000011100001100111110110011111010111011100100101000110110011000011001111110010110001100000011011001010011010100010101011001011110011100011000110110011111101001011001110001101110010100010011111100110000001011010010110100101100001011000010110000101010001011000010101100101100001011000010110100101101001011100010111000101110001011100010111100101110001011100010111000110000001011110011000000110000001011110010111100101110001011100010111000101110001011100010111100101110001011010010111000101101001011000010110000101100001010100010101000101100001011000010111000101110001011100010110100101101001011100011100001010010011011101001000010101011101000011001010110001111100000000111000001101010011001010100111100101111100010111001111110011100100110111001101110011010100110101001100110011000100110001001011110010100100100111001010010010000010101110011100010000000100011011000101110001010,
	960'b001000100011011111101100111110101110110000110001000111000010001000100011001001000010001100100000001101011110110011111010111011010011110000100110001011100100001001011000010101100010100100110101010011010101000001010111011000010111110110000100100010011001010010100101101010001010011010100010101000001010001010100100101001101010011110100111101010101010110010101110101100001011001010110100101101001011010110111000101110011011100110111011101110111011110010111101101110111011101110111100101111001011101110111001101110011011101010111001101110001011100010110101101101001011010110110010101100011011000010101111101011001010111010101101101010111010101010101000101001101010001110100010101000101010011110101010101001111001111010001110100011011001001010000110011010110110000101011101010111110011000100110010100110001010000110011111100111101001110110011101100111001001101010011010100110001001011110010101100101001001010010010011011010010011000001110101100011011000110010001011,
	960'b001000100011010111101100111110101110110101000011001100010011010100110101001101010011010000110100010001011110111011111010111011000011100100100111001011010011010100111101010011010011111000101000001010010100001001011100010111110110001001100110011010000111000010000100100100011001011010010111100101101001011010010111100100111001000110001110100010011000100110001001100010101000110010001101100100101001010010011011101000011010010110101011101011001011000010110000101100011011000110110100101100111011001110110001101100001011000010101100101010101010010110011110100110101001100010010001100011101000101110000111100001001000011110000110100010001000110010010000100100101001010010010100100101011001011010010111100100011000001001101100011001110110011101100000011001010101000100101110001101101001000010011100101000101010001010100001101000001001111110011110100111011001110010011011100110101001100110011000100101111001011010010101011110000010111001100101100011101000111010001100,
	960'b001101010100000111101101111101111111101111101101111010111110110011101100111011001110110011101100111011011111101111110111111011000011100100101001001100100011001100110111010000110011111000111101001001100010010100110001010011010110000101100000011000010110011101110010011101010111011101111010011110110111101001111001011100110110111001101010011001110110011101100111011010000110101101101101011100110111011001111100100000011000011010001110100100001001001110011000100110101001101110011100100110001001011110010101100101001001001010001110100011011000100110000000011110010111011001110001011010110110100101100111011001100110100101101001011010100110111101110001011100110111011101110111011110000111011101110110011101010110111101100000010101110101111001100100001111000010110100110110100100111010100010101000101001011010010010100011101000011010000110011111100111101001110110011100100110101001101010011001100110001001011010010110100000110011000101010001100011101000111110001110,
	960'b001010000011101111101111111110101111011111111010111110101111101011111010111110101111101011111010111110101111011111111001111011110011101100101000001100000010111100110000001101110011101000111110010000010011101100101011001010010010010000110000010100000111100110011010100101101001000010010000100100011000111110010000100011101000110010001100100010111000110010001100100010101000101110001100100011011000111010010010100100111001010110011010100111011001111110100001101000111010010010100100101000101010001110100010101000001001111010011001100110011001100010010101100101001001001010010001100100001000111110001111100011111001001010010011100101001001011110010111100101101001100010011000100110001001011010010111100111111010001101111010010010000010101000100011001110011001011010100011101010101010100110101000101001111010010110100100101000111010001010100001101000001001111110011110100111011001110010011011100110101001100010010111100011000011110001000000100011001001001010010000,
	960'b001010000011011111011101111011011110110011101101111011011110110111101101111011011110110011101101111011011110110111110000111000000011101100101100001011010010101100110000001100110011100000111011001111000011111100111110001011110010011100100100001000110010111101011010011100110111111010000011100001001000001010000011100001001000011110000010100000000111111101111110011111011000000001111101011111100111111010000010100001011000011010001101100011101001000010010011100101101001011110010111100110001001010110010011100100011000110110001011100010101000011110000110100001011000001110000001100000001000000001111111100000001000000110000011100001001000010010000100100001111000000110000010100000111000010001111110011100110101101100101010001010010001111000110011100110111011000110110000101011101010110010101100101010101010100110100111101001011010001010100010101001011010000110100000100111111001111010011101100111001001101010011010100101010100110000110011100001101001010010010011,
	960'b001101100010110100110110001110100011110000111110001111110011111100111110001111100011110101000100010000110100100101010110010011100011000100110000001010010010110100110010001110000101001101010011010000000100000101001110010011010011000100101111001010110010100100101000001010100011001001001111010001000010111100110000010001000100111000110011001011110011001000110011001110110100111000111000001100110011010000110110001101000011101101010000001110110011011000111000001110100011100100111111010110000011111100111000001110000011100000111001001111110100110000111110001101100011011100110110001101010011100101001001001110110011010000110110001110000011110101001101010101000011011000101110001111110101011100111011001100110010111000111010100100010100100010011100101100101011000110110000101100001010111110101111101011101010101010100011101000011010001110100011101000111010001110100011101000111010001010100001101000001001111110011111100111110110010100101101011111111001101010011001,
	960'b010001010010101000100110001010000010101000101100001011000010111000101111001011010010111000110111010000010011110000111101001111100011010000110010001010010010111000110000001110010110100101101111010010100100110001100100011000100100010101000011010010100100111101010101010101110101101101011101010110110101001001001001010000010100111001010110011011011000110110010100100100001001101010011001100100111010000010011101100100001001000110010101100101001001010110011000100110111001110010011111101000111010010010101000101010111010111010101111101011111010111010101010101001111010011010100111101001111010100110101011101010011010001110100010101000111010001110101000101011111010001001001011011010001011011010111000101110001011101110111101110001101011111111001001110010001100100111001001110010011100100011001001110010001100011011000011110000111100010011000101110001101100010111000100110000111100001011000000110000001011111111000000101111111000101000101100100001011011111010111011,
	960'b001111010011010100110111001101110011011000110101001101100011101100111100001111000011111101001010010100010100010001000000010001000100001001000001001110000011011000111000010000000100111101010100010010000100110001011000010101100100111001001111010100000101001101010111010110110110000001100101011011110111001001101100011010010111111010010001101011001100000111000010101110101011011110110100101100101100010111001011110010011100110111001101110011011101000011010101110101111101010111011000110110011101111011100001111001001110010011100000110111101101110111011111110111101101111111100000111000111110010011100100111010001110011011100101111001111110011111100111111011001110010101101111011101111110110011110100111100101111001111110011111100011111000111110000111011111111000011101111111011101110110111101100111011001110110011101010111010101110100011101000111001101110010111100010111000011110000111100000110111111101111111011111110111111011000000110001011111001101011011010110,
	960'b001111100100001001000100010000110100010001000101010001100100011101000110010001110100101001001100010011000100111001010000010100000101001001001111010001110100101001010100010101100101001101010111010101110101011101100001011001100110010101101000011100000111100001111100100001101001110010100010101011011011010010110011101100101011010110111000110000011100010010111110101110011011011010110101101110101100010111001011110011101100110111000110110010001101000011010100110101111101100011011111111001101110110011101111111101011111010011101111111011001110110111110000111011111110111111101010111100011111001011110011111100111111001111110011111011111110111011101000111010011110010001111110011001101110010011101010111010001110100011100111111010011110100111101001111010111110110011101100111010111110110011101100111010111110101111101011111010111110101011101001111010001110100011101000111010011110100011100111111001111110011011100110111010001100011100111101011001011101100011100000,
	960'b010011000101000101010110010110110101110101011111010111110101110101011011010111010101110101011010010101110101101001011111010111100101111101100001010111110110001101110001011110010111100001110110011101010111100101111110100001111001010010011100101011001011010110110101101101001011111111000111110010011100101011001011110011011101000011010001110100111101010111010001110011111100111011010001110101011101001111010101110101101011110010101000110000001101011011011110111000011110001111101000111010101110110111110000111101111111100011110010111100001111000011101111111100001111001011110001111100101111001011110010111100101111001011110001111001011110010011100010111000001101111010001111010101111101011111100001110111011101110011011001110110111101101011010110110101011100111111001000110010001100100011001010110010011100010111001011110011011100110011001101110010011100011011000110110001101100011111001001110010111100110111001110110100001011101101000110010101001101000111011101,
	960'b011010100110111001110010011110110111111110000111100100001000111010001101100011111000111110001110100011101001001010010100100101001001010010010100100101011001001110010110100111001001111110011111100111111010001110100111101011011011010110111011110001001100100111001001110010011100101011001010110011011100110111001101110011111101000111010100110110001101011111010110110101001101000111001011110001111010110110100100101001101001111010110011110011011101101111100011111001111110011011100101111001101110100111101101111101011111100011110001111100001110100111000011110010101101010111101000111100111111000111110000111100001111000011110000111011111111000011110001111100101111001110101111010100101101101011110100111100011111000111110000111100001111000011101111110111111010000110010111101010101010010110010100100101001010001110100011101000001010111110101010101001001010000110101100101011001010101110101011101010001010010010100111101010001010000101001110001111101010011110111010,
	960'b100101101001011010011000100111101010000010101000101100111010111110110001101101101011100010111001101110011011101010111100101111011011110110111100101110111011101010111001101110101011101110111110110000001100000111000011110001011100011111001000110010111100110111001101110011101100110111001011110010011100011111000110110010001100101111001001110010011100101011001000110001001100001010111100101111001011110010111101101110001010111110101101101010111010101010101010101011111011000110110010101101001011111111001100110100001101011011010001110011111101001011001001110100001101101011100111111011111110111011101100111010111110101011101010111010111110101111101010111010101110101010110101010010001100100011101011111001101110010111100110111001101110000011010011101100000111011001100101011001100110000101011001010110000101101001011000010110100110001101011111010111010101110101101100011100110111000001101010011000110110010101110100011110111000010001001110001011111000011110011111,
	960'b110001011100010111000100110001001100010011000101110001111100011011000111110010001100011111000111110001111100011011000110110001011100010011000100110001011100011011000101110001101100100011001000110001111100011111001001110010111100110111001101110011011100111111010001110100001101000011001010110001001100001111000100110001011100100110111111101110001011100111000000110000111100010111000011110000111100011111001001110001111100001111000010110000001011100010100011100101101000111110000110011111111000011010001101100010101000110010001001100010001001001110010101100101111010001010101110101111011100011011001000110000101100001011000110110010101100011111000010101111101011110110011011001110011001100010111110101101011011010110111000101100101010100010100000100101011000111110001011100010101000011010000100011110100111001001101011011000110101111101011011010110110101100101010110010101110101011101010111010110000101100101011000010101110101011100111110001001100101010001100110,
	960'b110001001100011011001010110011101100111111010000110100011101000111010000110011111100110011001011110010101100100011001010110011001100110011001100110011001100101111001010110010111100101111001001110001111100010111000010110000101100011011000110110000111011111110111000101011101010101010101000101010001010110110101101101101101100011011000110110000001011101011000111110011101100111111001101110011011100111011010000110100001100111011001110110011111101000011001000110000101100001010111101101100001010100010101000101010101010001010011011100101111000100001110001011011000111001101110011011110000111110110000101100010101000101110010000100100111001001010010010100100101001010001111101001100000111001110001111100000100111111101111110011111110111111001111011011101000111010001111011100000110111111010000010100010001000110010000010011100000111000001101111011101010111111101111111100000011000000001111111100000011000100110001111100001100111101001010110001001010101101101110110,
	960'b110001111100011111001000110010011100101011001011110011011100111011000011101100001010011110100110101000101010000110101100101100111011100010111010101110101011011110111000110001001100110111001011101111101010101110100011101010101011010110110111101100111010111110101010101000011001101110100001101100011100011111000110110011111101001111010011110010111100000111010010110111101101111011011010110110101101101111011100110110111101110111011110110111101110000011011111110111011101110111100001111000001101110011011011111001001110000011011000110100101100000010011001011111000111001101101101011010100110101001101100011100010111001101110011011100100111000101110100011100110110111101011101001010110100101101100100010111000101101101011011010110010101100001011010010110000101010101010011010101010101010101010110010110010101110001011001010101100101010101010110010110010101111001100001011000010110000101100110011011000111010101110110011100000110111101011001001001010100101101100111,
	960'b110010011100101011001011110011001100110111001101110011001100101110111100100111001000000001101101011001000101111001100010011010110111100110001001100100001000101110001100101011001100000010111111101011111001100010010111101010001010110110101111101011011010110010100111100110101000101110010101101010011100100011001011110111001101111111011110110101001100101111011001111001001110011011100100111001011110011111100110111001101110101011101100111010011110101111101011111010101110100011100111111001111110011011100101111011111110110111100100111000001101011111001001101110001010110110011101100010101000001101111100011110000111000001101011011010100110100101101000011001100101111101010011001011000011110101011100010101110101010001010011010100010101000001001101010010110100100101000110010001100100100101001011010011100100111001001100010010110100101101001100010011010100111101010010010011110100101101001011010011000100111101010011010100110101010001001001001001000011101001010100,
	960'b110001011100011111001010110011011100111011001110110011111100111111001111110011001100001110101001100011000110110001011101010111100110110010000001100011001000101001111111100010111001000010010001100011011000100110001100100100101001001110010110100110101001111110100010101000011001110010100000101110011101101111011011111000101110010011100100110111001101001011011111111010001110100111101000111001101110011111101000111010001110100011101001111010001110100011100110111001101110011111100101111001001110010011100100111011101110111111100111111000101101100111010100110100001100110011000111101110111011001010100100100101101000011110000000011101110111000001101101011001110101111001010101001100000011011001011001010101110101001001010010010011110100110101001010010001100100010001000011010000110100010001000101010001100100011101000111010010000100100001001001010011000100101101001000010001110100011101000111010001110100100001001010010010110100110101000111001001010011010101001111,
	960'b101111001011110010111110110000011100001111000101110001111100100011001001110010101100100110111100101010111001101110001110100001111000000010000110100100011001000110010011100100001000110010001000011111110111001101101010011011000111110110001011100011101000111010001111100100111001000110010101101001011011101110111101101101101011011011000101110010011100001111010000110111011101111011011001110110101101110111011110111000011110001111100100111001101110011111100111111001101110011111100111111001101110011011100100111011011111000111101100111010011110010011100011111000011110000111100000110101011100100111000100101111111011001110100110100110011001000110001011100001000111101101110000010000010011011001100110011000100101100101011000010110000101001101001110010010100100011001000101010001110100011101000110010001000100000101000010010000110100001101001010010011010100011101000001010000100100001101000100010001000100010101000111010001110100100001000011001000010011000001001011,
	960'b101110111011101010111001101110011011100010111001101110101011101110111100101111101011111111000000110000001100000111000001110000011011111110111110101111101011101010110010101001111001111010010101100100001000101010000011100001011001000110010111100101011000111010001000100000010111011001110000011100100111100001111001011101100111011001111100100001011000100110010111100110101001100110011001101110011011101010110101110000101100110011010010110111001110001111100011111000111110001111100001111000001110010111101010111100001111000111101100111010101110011111100111111001101110010011100010110111011101011011010111110111001101100011001010110000011100010011000011101110011010111010100010011000100011110010000111100011001000011001111100011100110110101101100010010110010101000101001110010100010101000101010011010011100100101001001011010011000100011101000110010001010100001001000000010000110100001001000000010000010100000101000001010000100100001100111110001000010010111101001011,
	960'b101110101011101010111011101110111011101010111011101110101011101110111100101111011011110010111101101110111011110010111110101111111100000111000011110001011100100011001000110010001100011011000010101111101011100010110000101001101010001110100000100110111001101010011111101000111010001010011011100110001001001010001100100010011000001001110110011011100110100001011111010110110110001001110100100000100111010101110111100010011001111110100110101101101100000111001111110101111101001011001001110011111101111011100111111100001111001011101101111011001110100111100110111001001110000111100001111000011101111111011101110111001101010011001101110001101100011011001110110011101100101111000111100001010100010010110111110011011100011110111101101100111010111010100011100100011000101010000011011111010111101101110110011011110110110001101010011001110101111101011000010100110101000101001111010011000100011101000100010000110100001101000010010000110100001100111100001000010010111101001010,
	960'b101110111011101010111011101110111011101110111100101111101011111111000000110000001100000110111111101111011011111010111110101111111100000111000011110001001100011111001000110010101100101111001100110011101101000011010011110101101101011111010010101111101010011110100000101000101010001110101011101011111011011010111000101111011011111010111011101101101010111010100000100100101000101010001110100010110111001001100111011001110110100101101000011100100111111010001110101000001010000010011110101011101011110111001110111000111110100011100011111001001110001111011110110110111101011011010001110100111101010111010110110110111101111011011100110110111101110011011101110110011101001111010001100110100100010010111011110100111100101111000111110010011100110111000101101110111011100010111000101011111010001010011001100101111001011110001101011111010111011101111101100000010111111001111011011100100110100101100011010110100101000101001110010010000100010100111100001000010010111001001010,
	960'b101110101011101010111011101111011011111010111110101111111100000011000010110000101100001111000011110000111100010011000100110001011100010111000110110001101100100011001001110010101100101111001101110011011100111011010000110100111101100011011011110111001101101011010101110100001100100011000100101110111011111110111110101110101011111111000111110011101101100011011111111000101101110011010110110011111100001010110011101001101001011110000110011101110111000101101100011011000111000001110101100000111001010010100001101011001011101011000010110000111100011011001100110100111100111011000001110000111100011011001000110011011101011111011101111000001110000111011110110110101101011011011001101011010100010010110010110101001100111011001110110101001101011011010000110011001100011111000001101111111011100110110100101011101010101010100111101000101001111010011111101000111010000010011011100110001001011110010001100001110111111001110101011011000110100001011001001001010011010001100010,
	960'b101011001011010010110111101101001011010110110111101101111011011110111101101111111011111111000000110000011100001011000011110000111100001111000100110000111100010011000111110010011100101111001100110011001100110111001110110100001101001011010100110101101101100011011000110110101101111011100001111000101110001011100010110111001101100111010101110101011101100011011110111011101111010011110000111011111110110011101001111000111101110011010010110001011011100110100110100011001000001110000101100001101000110010001011100000001000000110001100100100101000111110010001100110001010100010111101101110001010101010101100101011011010111110101110101101001100100011010011110010011011011010111111101010000011111110011101110010111100010011000001110001101100101011001010110010001100001110111111110001001100110011001000110001011100010011000000101111011011101010110101101100001011000010101101101010111010101110101010101010001010001010100000100111011001100001111100001010100011110101111101,
	960'b101001001010101110101010100110011001111010100111101010111011001010110101101101101011010110110111101110111011111011000001110000101100001111000011110000111100010011000101110001111100100011001001110010111100110111001111110100011101001111010101110101101101100011011000110110101101110011011111111000111110011011101000111010101110101011101001111010001110011011101001111100001111010011110011111100111111001011110011111100111111001011110001111100001110111011101011111001011101110011010000110000011011101010110010100111111001010010010000100100001000100101110111011100010111110010000010100000000111101101111100011110010111010001111000100000001001011010100100101011101001111110011101100011000011100010001001101111011011011010110000101101011011111011000100110001011100010011001010110011111101001011001110110010101100100111000011101111011011100010110110101101111011111010111111101110111011101010110110101100111010110110101011101010101010100110001011001011100100011110001110,
	960'b101010111010100110101001101010101010110010101101101010101010111110110100101100111010111110101111101101011011100010111011101111001011110110111101101111011011111011000001110000111100010111000111110011001101000011010100110101111101100011011001110110111101111011100000111000011110001111100100111001101110100011101010111010111110110011101101111011011110110111101110111011111111000011110000111011111110111011101110111011111110111111110000111011111110111111110000111011111110111111101011111000111101110011011000110101011101000011001011110001111011110110011101100011101000000101110001011010010110011001100001010111010110000101101010011110111000110001111111011111011000000010000011011110110011011101101000100101001000101110000010100010101001111110110000101110001011111011000000101101101011010010110110101011011010110110110111101111011011101010111001101111001011110010111000101110011011101110110110101101011011011110110110101101001011000110001110001011010100111010010111,
	960'b101010111010010110011111101001001010100110101100101010111010111010110100101101101011011110111001101110011011100110111001101110011011100110111011101110111011101110111100101111011011111111000001110001101100111011010100110101111101100111011001110110111101111111100011111001101110100011101001111010101110110011101101111011101111000011110001111100101111001111110011111100101111001011110010111100111111001011110000111011011110110011101011111010011110100111101000111010001110011111100111111001001101110011010110110101101101010111010110110101001101001011001110110010101100001010110110100111101000101001111001011100000110111101100101011001010110110001101001011010100110111101111000011100110011010101010011011111100111110101111100100000101000010110000110100010111000110110010100101000011010111110101111101001101010010010101000101011111011001110110101101110101011110010110101101100011010111010101110101011101011000110110010101100011011000010001010001010000100110110100001,
};
parameter [0:85][959:0] g_picture = {
	960'b011110101000010010000101100001011000001001110101010111110100101100111011010001110111100110000110100010001000100010001001100010101000101110001100100011011000110110001110100011111000111110001111100100001001000010010001100100011001000110010010100100101001001010001101100000111000001010001011100101001001011110011001100111001001011110001111100011001000110110001100100100111001100010011101100111111001110010011111101001011010110110110010101011111010100110101010101100101100000011000101110000011011111010111100101110101011100010110110101100111011000110110000101011011010101010101000101001101010010010100010101000001001111010011101100110111001101010011000100110001001011010010101100101001001001110010011100100101001000010010000100011111000111010001110100011001000101110001011100010101000100110001000100010001000011110000110100001101000010110000100100000111000001110000011100000101000000110000000100000001000000001111111011111100111111001111110011111010111111001111101,
	960'b010001000101111010001000100011101000110010000011011100110101111001001010010100000111110110001101100011111001000010010000100100011000101110001011100011001000110110001110100011101000111110010000100100001001000010010000100100011001000110010001100100101000111010000010011111010111111010000001100001111001000110010110100110001001011110010011100100111001001010001110100101001001110010100110101010101010100110101100101101001011100110111111101110111011011010111000110000001100100011001001110001111100010011000010110000001011111010111100101110011011010010110001101011101010110010101001101010001010010110100010101000011001111010011101100110111001100110011000100101111001011010010101100100111001001110010010100100001001000010001111100011111000111010001101100011001000101110001010100010101000100010000111100001111000011010000110100001011000011010001100100010111000101110001010100010101000100110001001100010011000100010001000100001111000011110000111100001010111111101111101,
	960'b001111100100010011001111111000001101111011011110110111011101101111011001110110011101110111011111110111111101111111011111110101101001000010001010100011001000110110001110100011101000111110010000100100001001000110010001100100011001000110010001100011111000011110000000011111100111111110000000100001011000111110010101100110001001110110011101100111001001111010011010100110001001100110011100101000001010110010110100101110001011111111011110111000111110001011100011111000111110010011100100111001001110001111100011111000111110001111100011110111011011100110110010101100001010110110101011101010011010011110100100101000011001111110011101100110111001101010011000100101111001011010010101100100111001001010010001100100001000111110001111100011101000110110001101100010111000101010001010100010011000100010000111100001101000011010000110100001001000110011010101110111111101111011011110110111101101111011011110110111101101111011011110110111101101111011011111110101011000010101111101,
	960'b010011110101010011011010111110011111100011111010111110101111101011111011111110111111101011111001111110011111100011111000110111111001000110001010100010111000110110001110100011101000111110010000100100001001000010010000100100001001000010010000100011101000110010001010100001111000100010001100100011111001011110011011100111101001111110100001101000101010010110100110100111111001110110100000101000011010100110110100101110011011111111100011111110001111011111110111111101111111011111110111111101111111011111110111111101111111011111111000111000101011101010110100101100011010111010101100101010101010011110100100101000101010000010011110100111001001101010011001100101111001011010010100100100101001000110010001100100001000111110001111100011011000110110001100100010111000101010001001100010001000011110000101100001001000001110000100100000111000101111011111111110011111100011111001111110011111100111111001111110011111100111111001111110011111100011111001110111111000011001111101,
	960'b010111000101101111011010111110011110011111011001110110001101100111011000110101111101100011011011110111111110011111111000110111111001000010001010100010111000101110001100100011101000111110010000100100001001000010010001100100001001000110010001100100011001001010010010100100111001010010010110100101111001101010011100100111101001111110100000101000101010010010100111101001111010100010101100101011011010111010110101101110011100000011100011111101111110100011100100111001001110010011100100111001001110010011100100111001001110100011110111111000111011101110110100101100101010111110101100101010111010100010100100101000011001111110011101100111001001101010011001100101111001011010010100100100111001000110010001100100001000111110001110100011011000110110001100100010111000101010001001100001111000011110000011011111000111101110000001100000111000101111011110111110001110011111011111110111101101111011011101110111011101111011011110110111101110011111111000110111101000011001111101,
	960'b011001100110010011011010111110111101100101001100010001000100101101000000001110000100001001100001100001111101111011111001110111000111011101111000011110000111000001101111011101010111110010000111100100001001000110010010100100101001001010010010100100111001010010010101100101101001011010010111100110001001100110011011100111011001111010100000101000101010010010100111101010011010101110101110101100011011010010110101101110011100000011100011111101111110010011001010110010111101000111010110110101001100111111001011110010101110010011110111111000111011101110110100101100101010111110101100101010101010011010100100101000011001111110011110100111001001101110011001100110001001011010010100100100111001001010010001100100001000111110001110100011011000110110001100100010111000101010001000100001111000011010000011011111000111101101111110100000011000101111011110111110011101111110001111100001011000001001111011011111011000001110000000100001011101111011111001110111101000010101111010,
	960'b011011010110111011011100111110101101011100111001001010100010111100101001001000110010101000111010010101011101101011111010110110100101011101000000001111000100010001001001010011100101100001100001011111011000111010010000100100011001000110010010100100111001010010010101100101101001011010010111100110001001100110011011100111011001111010011111101000101010010010100110101010011010110010101110101100011011010010110101101110011100000011100011111101111110001111001000110101011110001111100101111000101101011111001000110001101110001111110111111000111011101110110100101100101010111010101100101010011010011010100100101000011001111110011110100111001001101110011001100110001001011110010100100101001001001010010000100100001001000010010000100011101000110110001100100011001000101010001000100010001000011010000100100000111000001010000010100000011000101011011110111110011101111010000011011101100111001001101111011100000111001101101111011110011101110111111001110111010111111101110010,
	960'b001110010101100111011011111110111101011000110001001001110010011000100001000111110010010100100110001110011101011111111011110110000011110100101011001101000100001001001111010101010110110001101100010111100111111110001111100100001001000010010010100100101001010010010101100101011001011010010110100110001001100110011011100111011001111010011111101000101010010010100110101010001010101110101101101100011011001110110101101110001011111111100011111101111110010011010000111001011110100111100111111001101110000111001101110001011110001111110111111000101011101010110011101100011010111010101100101010011010011010100011101000011001111110011110100111001001101110011010100110001001011110010101100101001001001110010010100100011001000110010000100011011000110010001100100010111000101010001000100010001000011110000111100001101000010110000001011111001000000111011101111110011101110101111101011100010111001001110001011100000111000001101110011110011101110111111001110111010111100101101110,
	960'b000110110011000011010111111111001101011000101100000111110010010000011100000111010010010000100010001101001101011111111011110101110011110100110110001111110101001001100100011010000111001110000100011110010111001110001011100100001001000010010001100100101001001110010100100101011001010110010110100110001001100010011001100111001001110110011111101000011010001110100101101010001010101010101101101100001011001010110100101101101011110111100011111101111110010011010110111010101110101011101000111001111110010111010000110001011110001111110111111000101011100110110011101100011010110110101010101001111010010110100011101000001001111110011110100111001001101010011010100110001001010110010110100101011001001010010001100011111000101110001000100010011000101110001100100010101000100010001000100010001000011010000101100001011000001101111111011101110111110011011101111110011101110101111011011100010111001001110010011100000110111101101110011101011101110111111001110111010111101001110001,
	960'b000110010010101011010110111111001101011000101100000101100001101100011011000111000001111100011101001100001101011011111011110110000011111100111100010010110110000001110110100000011000010010001010100011101000100110001101100100001001000010010001100100101001010010010101100101011001010110010110100110001001100010011001100110111001110010011110100111111010001010100100101001101010100110101011101011111011000110110011101101101011110111100011111101111110010011010101111010101110101111101001111010001110010111001111110001011110001111110111111000101011100110110010101011111010101110101000101001011010001110100001101000001001111110011100100110101001101010010101100010001000010010001110100011011000111010001110100010011000000001111000011110101000010010001010100000100111110010000001100001011000011010000100100000100111111101111000011100010111101111011101111110011101110101111011011100010111001001110001011100000111000001100100011000111101101011111010110111010111101101110001,
	960'b001100110011011111010111111111001101011000101000000101000001011100011010000111000001110100011011001100011101011111111011110110000100001001000000010111000111010010000011100010101000110010001110100011111001000010010000100100001001000110010001100100111001010010010100100101011001010110010110100101101001011110011000100110101001101010011100100111111010000110100100101001011010011110101010101011011011000110110011101101011011110011100011111101111110010011001101111000111110110111101100111010101110000011000111110001001110001111111000111000101011100010110000101011011010100110100111101001001010001010100000100111101001010010001110100100001001001110000011011101010111100101111101011101110111111010000110100000100111100001110011011101000111101010000001011101110111001101110101011110101000010010000010011110100111011001110011011100000111101011011101111110011101110101111011011100010111001101110010011100000101101101000010010101101101101011111010110111010111101101101111,
	960'b010110000101001011011001111110111101011000100110000100100001010100010111000110100001101000011001001011111101011111111011110110010100110001001011011011111000001110001011100011001000110110001110100011111000111110010000100100001001000010010001100100111001001110010011100101001001010010010101100101011001011010011000100110011001101010011011100111101010000110100011101001011010011010101001101011001010111110110001101100111011100111100010111101111110001111000110110011001101111111100110110111111100110011000001110000011110001111111000111000101011011010101110101011001010100010100101101000111010001010100000100100110111110001110111100000011000010101111001011101000111010001110011011100110111010101110111011101100111010001110011011101000111010101110110011101010111001101110011011101100111110101111100011101010111001001110010011100000111101011011101111110011101110101110110011011100111000001101111011001010011110100110110010100111101101011111010110111010111100001101100,
	960'b010000110100111011011001111110111101011100111011001001110010100100101101001011010010110000101011001111011101011111111011110110000100001001000010011001100111111010001001100011101000111010001110100011111000111110010000100100001001000110010010100100111001001110010011100101001001001110010101100101101001011110010111100110001001100110011011100111101010000010100010101000111010010010100110101010011010101110101110101100001011011011100010111110001110001111000101110001001100100111001100110010011100010111000001110000101110001111111000111000101011010010101011101010011010011010100100100110111001110010011101100001010111010101110100011110000111100001110101011101000111001101110011011101000111010001110011011101000111001101110100011101010111010101110101011101000111001101110101011101100111011001110101011100110111000101110001011100000111101011011101111110101101110001110011011101000111100001110111011001000100010101000101011000001101101111111010110111000111000001100110,
	960'b000110010010110111010110111110101110011111011000110101101101011011010110110101101101011011010110110110001110011111111010110101110011101100110011010000010100101101100000011110101000011010001011100011111000111110010000100100011001000110010010100101001001001010001111100010011000010010001110100101011001011010010110100101111001100010011010100111001001111010011111101000001010001010100100101001111010100110101100101011011011010011100010111110001110100011100011111000111110001111100011111000111110001111100011111000111110100011110111111000101011000110101000101001101010011010011011100000101000110110010101011111100111011001110110011101000111001101110100011101010111010101110011011101000111010001110100011101000111010001110101011101010111010001110100011101000111011001111000011101100111011001110101011100110111001001110010011100100111110011011101111110011110011111011100110111001101110111011101110110111101100011011000110110101110011111111001110110110110110001100100,
	960'b000110110010111011011000111111001111100111111011111111001111110011111100111111001111110011111100111110111111100111111011110110010011111100111001010010010100100001001000010110010110110001111001100001111000110110001110100011101000111010001110100100001000111010000011011110010111100010000010100100111001011010010111100101111001100110011011100111011001111110011111101000001010001010100011101001101010100010101010101010111011001011100010111110001111011111111000111110001111100011111000111110001111100011111000111110001111011111111000111000101010111010100110101000111001101110001011011101111000000010001011100000000111100101110110011101010111010001110100011110110111110101110111011101010111011101110100011101010111010001110100011101010111010001110100011101010111100001110111011101010111010101110101011101000111010001110100011101000111111011011111111110101111100111111010111110101111101011111010111110111111101111111011111110111111100111111010110111010110101101100010,
	960'b001110110100110111001100110110011101011111010111110101111101011011010110110101101101011011010110110101111101011111011001110010100100100000111100001111110011111001000100010100010110001101110011011101011000010010001100100010111000011010000100100010011000110001111111011101010111010001111011100011101001000010010100100101111001100010011010100111011001111010011110100111111010000110100010101001001010011010101000101010011010111111011100111000101110001011100010111000101110001011100010111000101110001011100010111000101110000111100010110110111010110010100001100101011000001001111001011110011000010110001101100010101000000101111011011110010111011001111000011111010111101101110101011101000111010101110100011101000111010001110101011101010111010001110100011101000111011001110101011100110111010001110100011100110110110001100001010110010110001011001011110110101101101011011010110110011101100011011001110110001101011111011000110110001101100011011010110100000110110101011111,
	960'b010111100101100101001101001100110010111100110111001100110010101000100101001001100010011000101111001100100011000100110111001111110100000101001111010011010100010000111111010000000101000001110101100000001000000110001001100010101000000001111010011111001000000001111001011101110111011101110100011110001000010110001011100100101001100010011000100110101001101110011100100111011001111110100001101000101010001110100101101001101010011110101101101011101010111110110000101100011011001010110011101100101011001010110001101011111010110010101011101010101010000110010000100000000111101101111010100000101000111110010100100100111000110010000101100000000111110101111100011110000111010001110011011100110111010001110100011101010111010101110101011101010111010001110100011101000111010001110011011100110111001001110011011010110101100001000111001110010011001000111011010000110101001101010111010010110011111001000011001111010011101001000000010000110100010101010000011001010110000101100011,
	960'b001101010010011000011010000101110001011100011010000101100001010000010011000100110001010100011110001010000010011000101001001010110010100100110001010001010101001101011001010101010100011101100000100000111000011110001001100010101000011110000001011110010111001001101010011011100111011101100011011000100111100101110101100010011001100010011001100110101001101110011100100111001001111010011111101000001010000110100010101000111010010010100100101001101010011110101000101010011010101110101011101010101010101010101000101001011001111110011010100110101000110110000010011111010111110101111111100001011000111110010010100100011001000010001010100001100111110101110001011011100111000101110011011101000111001101110000011100100111010101110101011101010111010001110100011101010111010101110011011100110111001001110010011011010110100101100011010110100100101100110111001001100010001000101101001101000010101100100110001001010010010100101010001011000011001001000101010101000101110001011111,
	960'b000110100001101000011101001000110010010000100001000110100001100000010111000101110001111000100101001100110100011001000100010001110011101000110001001101000100010001010101011001110101111001001001011010101000001010000101100010001000011010000011011101100110100001100000010111100110101001011011010101110110001001110011100011101001011110011001100101111001011110011010100110011001100010011110100111101001110010011110101000011010001010100011101001001001111110010111100111101010011110101001101010011010100010100110101000101001101110010100100101011001000010001000100001011000011010000011100001001000100010001000100010001000100110001001100001110111110001100110010011000101010101101000011100000110010001010111011000110111010101110110011101010111010101110101011101010111010001110011011100110111001001110010011100100111001001110001011010010101001101000011001101010010010100011100001000000010001000011111000111110010010000101001001010010011001101000100010011100101000001001010,
	960'b001000100010011100110000001110010010100100011100000110100001100000011000000110000010100000111101001011000011100001000011010010110101011001001000001101110011100001001100011000000110110001011010010100110110110001111011100000001000000101111010011100110110111001100011010101010100111101001100010010000101000101100011011100111000011110010100100011101000110110001111100000111000000010010100100101111000011110000110100110001010000110100001100110101000010001111000011111101001000010100010101001001010010010100011101000101010000010011110100111001001101010010101100100011001000010001011100001011000010010000010100000000111111110000011100001000111110001100111010001010011010100111111010100110100001001000010011000110111010101101100011011100111010001110100011100010111001001110011011100110111001001110010011100100111000101110000011001110101111101010101010010000011001000100010000110110001100100011000000110110001111100100100001001100011001101000100010000010011001000101100,
	960'b001110100100011001001001010001010010010000011001000110100001100100011001000110000010110101011000010000000010101001000010010001010101001001011100010010010011010100111110010111000111000001110100011011000110100001110000011101010111011101110101011100100110110101100001010101100100100001000001010000010100100101010111011001000111011110001010100010011000011001111101011101100111010001111101100000010111110010000101100101101001111110011110100010110111010101110010011100100111100110001111100110111010000010011111100110111001101110011101100111011001101010010111100101001001001010010000100010111000100010000001011010110101110101101001011110110111111001110000010100110011001000101010001101010011010000111110010110010101111001010001011001110110111001100011010111000110011001110000011100110111001001110010011100010111000101110010011011110110111101101011010111100100110000111000001000110001101000011000000110000001101000011101001000010010100100101001001000100010000100100111,
	960'b010101100110000101010110001101110001110000011010000111000001110100011101000111000011011101100001010100000010100000101101010010000100101101010110011000010100100000110110010100110111011001111010011101100111001101101110011100010111000001110000011100000110101101100000010100110100010100111101001111010100010101010111011101111000001010000101100001101000001001110011011100100111000101110010011101111000100010011000100110111001001110010010011111110111001101110010011101000111011001111001100001111001010110001001011111110111111110001010100110101001100110010110100100111001000110001110100010111000100110000110011110110110001101010000010101010110101101101111010101100011001100100111001010000010110000110100010001000100011101001100010110000100101101001001010110000110101101110011011100110111001001110010011100010111000101110001011100000110111101101101011010000101100101000010001011100010000000011001000110000001100000100010001010000001110100011100001000100010100000110000,
	960'b011011000110100001000010000111110001101000100000001001000001111100011110001010000101011001101001010110100011100100100100001100000101000101010100011000110110011001000110010010010111010001111100011101010111000001110000011100100111000101110000011100000110111001100110010100110100101000111101001110010100010101001110011001110111100101111111100001010111100101101111011011110110111101110010011110101000100110010000100010010111100101111000011101000111000101110010011101110111010101110010011101100111110001110101011100100111001001111101100101011001011110010100100100101000111110001101100011001000100110000111100001100111110101100110010101010100111101011010010101110011001100100011001001010010101100101110001101010100001001000010001100110011011101010010011010110111011101110100011100110111001101110010011100100111000101110000011100000110111001101010011000000101011001001000001110010010011100011110000110100001110000110100001010010001110000100101001101110011111000111110,
	960'b011100000101010000100101000110010001111000101000001100100010000100011101001111010110101001101110011001110101011000111000001000000011011101011011010111100111001001100110010011110110101001110111011100000110110101101101011011100111000001110000011100100111000101101010010101000100010100111010001101100100000001010010010111010110100101101100011011110110101001101001011010000110100001101011011101010111110101110101011100100111100001111001011110010111101101111101100000000111111101111110011111110111111101111110011111010111110110000001100100111001100110010101100011001000001110000000011111110111110101111100011111000111101101110000011001010101101101001000010001000011011000100101001001100010011100101001001100010011100100101011001011010100000001011010011011000111010101110011011100110111001101110010011100100111000101110000011100000110111001101000010110010100110001000010001110100011000000100100000111100001110100101000000111100010000000101011001100100011011100111011,
	960'b010100000010111000011010000111100010100000110000001111000010011000100001010101000111000101110001011100000110110001010000001001110010001101000001010111110110111101110110011001010110000001101101011011000110110001101101011011100111000001101110011011000110110001011110001101110011000000110001001011110010110100110000001100010011000000110000001100000011000000101111001011100010111100101110001011100010110100101100010010101001001010110011101111101100100111010011110111101110010011100110111001111110011011100011110111011101000111001000101111101011011010011010010101000010111000101100001010110010101100101011001011010010111100101111001011110010111000101100001011010010101100101001001010000010100100101011001101000100010100101100001110000100101101100001011100000111001101110100011100110111001001110010011100100111000101110000011011110110110101100100010100010011110100110001001010110010001000011001000101010001011000010111000110010010001000101000001100010011110001000010,
	960'b001100000001111100011101001010010011100101000001010000000010010100100111011000010111000101110001011100100110111001100001001110100010001000101010010011110110100001110011011100010110010001101010011010110110101101101101011011010110011101010100001110100011011000111010001101110011011100111000001110010011011100110111001100010010111100101100001011000010110000101011001010010010100100101001001010010010100100101000001010010100001010000101100101001001100010011100101000101010001110100100101001011010010010100011101000011001110010011000100100111000010101000011001010010010100100101010001010010010100100101000001010100010101100101011001010100010110000101100001011100010111100101111001100000011000000110010001100010010111100101111010001100100101101001111010110010110011001101111011100010111000101110100011101000111000101101111011011000101101000111101001011010010011100100110001000110001110000010110000101000001010100010101000101110001100100011110001011110100011001001101,
	960'b001000010001111100101000001110100100101001010101010010100010010100111100011011000111000101110000011100010111000001101000010011110010101100101000001111000110001001101110011100010110011001101000011010110110101101101000011000110011011100111000001111110100001101001011010011000100111001001110010011000100100001001000010001100100011001000110010001100100010101000100010000110100000001000000010000000100000101000001010000010100000101000100010001010100011001000101010001010100010101000101010001010100010101000110010001110100011101000111010001110100010001000000010000100100001001000011010000110100001101000010010000110100001001000010010000100100001101000100010001000100010101000100010001010100001101000010010001000100010000111100001101010011000000110111001101000100010101011110011011110111010001110110011101010111000101101100010110010011011000101001001011010011101101000000001011000010001000011010000110010001100100011010001000000001110100011010000111010011001101001011,
	960'b001000100010100000110111010001110101100001100100010110100010110101010100011100000111000101110000011011110110111101101101011000110011110100101101001100110101001001101101011100000110101001101010011011010110010100111100001110110100100101100010100001011010001110111101101111011011011110101110101010111010101010101011101010011010100010100111101001111010011110100111101001111010100010101000101010011010100110101001101010101010100110101000101001111010011110100110101001011010010010100101101001011010010110100110101001101010011010100101101001101010010110100111101001111010011010100101101001001010010010100011101000111010001010100010101000101010000110100011101000111010001110100100101001101010101010110110101110111011010010001100011001110100101100111101001101000011000101000100011010100111011001110100011100100111000001011101001110110010110000110010010010010101110001001110001011000010001000011010000110010001100000100001001101000010101000100011000110110001110100100110,
	960'b001010110011100001000100010101100110000101101011011000000011100001100010011100010111000101110000011100000111000001101111011011010101000000110011001101010100100101101001011100000110111001101100011010100100100101000110010100111000011110101000101111001011100010010000011101110110101001100000010111110101111001011101010111100101111001011110010111010101110101011101010111100101110101011101010111010101110101011101010111100101110101011110010111010101110101011101010111100101110101011101010111100101110101011101010111010101110101011100010111000101110001011100010111000101110101011100010111000101110001011100010111000101110001011100010111000101110001011101010111100101110101011101010111110110000101110100100010011010001110111101101100011001001101101110010011100100010001000011011000110111001001110101011100110110010000111101001011110011011101001010011000000110010001001111001100010010000000011000000110000001100100100111010010100100011100111011001100000010001000011100,
	960'b001100110100011101010100011000110110101001101011010110010011110001101011011100110111000101110001011100010110111101101110011011000101111001000010001111100100111101100010011100000110110001011001011000000110110010011001101100100111110101011001010110010110100110000011100010101000111010001111100011101000110010001010100001101000010110000011011111110111111001111101011111100111110001111100011111010111110101111111011111111000000110000101100001111000100010001011100011101000111010001110100011101000101110001000100010001000010110000010100000010111111101111101011111000111111001111011011111000111110101111101100000001000000110000011100001101000100110001010100011001001000010001111100100011000111110001001100000110111011001011011010101100111010110100110101010001000000001101111011010010110110101110100011011000100010100110001001111010101001001100100011010110110011001011001001110100010011100011011000110100001110100101011010100100101111101011000010011100011010100100100,
	960'b001111100101101001100100011011000110111001101011010010000100001001101111011100110111000101110001011100000110111001101110011011010110101001010111010000110101100101101010011010110101110101101001011110011010010110111001100110000101101001100100011110111000101010010001100100001000111110001101100011011000110010001010100001101000010010000100100000010111111101111110011111100111110101111101011111110111111010000000100000011000001010000101100001111000100110001011100011011000110110001100100011001000101110001001100010011000010110000010100000101000000001111110011111010111111101111111011111110111111101111111100000101000001010000011100001101000100110001011100011001000111010001101100011111000110110001101100011001000100001111001011001010101010001100000101110101011100010010011100000100110100001110000010101100011100000111111010110000110100101110010011100100110111101011111001110010010001000011101000111010010001000110000010100010110100001101000010111110100111000111010,
	960'b010100000110011001101101011011010110111001100111001110000100111001101110011100000110111101101111011011110110111001101110011011010110111001100011010010110101100101101001010110100110011101111100101000001011000110000110010110100111101010001011100011111000110010000111100010011000110010001101100011011000111010001100100010011000100010000111100001101000010010000100100001001000010110000101100001011000010110000110100001101000011110001000100010101000101110001100100011011000111010001101100011001000110010001100100011001000100010000111100001111000010110000101100001001000011010000110100001101000010110000101100001111000011110000111100010011000110010001101100011101000111110001110100011111000110110001000100001011000010110001010100010000111110001101000011111011011010010110100100110000111110101100011010011010100001001011100011011100111011001111000011101100111001101011101001011110010000100100010001000010010100100111101010111010110110101101110011001100101110001001100,
	960'b010111010110101001101110011011100110111001011100001100000101110101101111011011100110111001101111011011110110111101101111011011110110111101101100010111010101111001000011011001110111011110010100011100100110010010000110100100101000100110001000100011101001000010000011011111010111110001111101011111010111110001111100011110110111100101111001011110000111011101111000011110000111100101111000011101110111100001111001011110010111100101111001011110010111101001111100011111000111110001111100011111000111110001111011011110110111101001111010011110010111100101111000011110000111100001111000011110000111100001111000011110000111100101111010011110100111110001111100011111010111111001111110011111100111110101111101011111111000011010001101100001111000011010001000100010000110100101101100101010011000101101111110011001010101001101110000011101110111100101111000011101110111010001011000001010100010011100110000001001010011000101001010011001100111000101110000011010110110000101011010,
	960'b011001100110110001101110011011110110110101001101001101010110100001110000011011110110111101101111011100000111000001110000011100000111000001101111011010100110001001000101011010101000101110100000011010001000101010011001100101001000101110010001100011001000000101111100011111000111101101111010011110100111100101111001011110010111100001111000011110000111011101110111011101100111100101111000011101100111011001110111011101110111011101111000011110000111100001111010011110010111101001111001011110010111100001111001011110010111100001111000011101110111100001110111011110000111100001110110011101110111011101110110011101100111011101111000011110000111101001111010011110100111101101111011011110110111101001111011011110100111101110000101100100001000110110001010100101111000110101100101011101011010010110000101011011010100000101100111011101110111100001111000011101110111001001001101001010010011010001000001001010100011101101010101011011000111000001110001011011110110100001100010,
	960'b011011010110110101101101011011100110100100111100010000110110110101110000011100000110111101101111011100000111000001110000011100000111000001110000011001100011101001000110100011101001011001101011100110011001100110010010100101001000010001111111011111100111110101111001011110000111100001111001011110000111100001111000011101100111011001110110011101110111100001111000011101100111100001111000011110000111100001111000011101110111011101111000011110000111100001111000011101100111100001111000011110000111011101110111011101110111011001111000011110000111100001111000011110000111011101111000011110000111100001111000011110000111011101110110011101110111100001111000011110000111100001111000011110000111100001111000011110000111100101111011011111011000000010001100100100001001011010011011100101011001111110110101100000110011111000110110011011010111011101110110011101010110110101000000001100000100101101011010001100000100001101100001011011110111000001110000011100000110110001100110,
	960'b011011010110110101101101011011010110000100110001010101000110111101110000011100000111000001110001011100010111000101110000011100000111001001101100001011100010111001001110100101000111100001111101100110011001010010010100100101101000000101111101011111010111110001111000011110000111100001111000011110000111100001111000011101100111011001110110011110000111100001110111011101110111100001110111011110000111011101111000011110000111100001110111011110000111100001110111011101110111011001111000011110000111100001110111011101100111100001110111011110000111100001111000011110000111011001111000011110000111011101111000011110000111100101111000011110000111100001110111011110000111011101111000011110000111100001111000011110000111100001111011011110110111111010000010100101001001001010011010100111010111001110101101101001000100000100101011001110110111000101110101011100110110011100111001001110110101111001101000001111000100101001101011011100000111000001110000011100000110111101101001,
	960'b011011000110110001101101011011000101000100110011011000110110111101101111011100000111000001110001011100010111000101110001011100010111000101100101001011000011110001101100011100011000110010011011100100101001100010001101100001000111111001111011011110100111100001111001011101110111100001111000011101110111100001110111011101110111011101111000011101100111011101110111011110010111100001111000011101110111100001111000011101110111100001111000011110000111100001111000011101110111011101110111011110000111100001110110011101100111011101110110011101110111100001110111011101100111100101110110011101110111011101110111011110000111011101110111011110000111100001111000011110000111010101110110011110000111100001111000011110000111100001111001011110100111110001111111100001101001011010010010100100101000111101110110101000110101000100101001001010110110100101110011011100100101100100110101010010000110011101101101010001010101000101110000011100100111000001110001011100000110111101101101,
	960'b011011000110110001101101011010100100001000111101011010110111000001101111011100000111000001110000011100010111000001110000011100010110101000101100001010010100110110000000011101101001101010011000100101001001001110000011011111110111110001111011011110010111100001111000011110000111100101111000011101110111011101110111011101110111100001110111011101110111011001110111011101110111011101110110011101110111100001110111011101100111011001110111011101110111011001110111011101100111011001110110011101100111011001110110011101100111011001110110011101100111011101110111011101100111011001111000011110000111011101110111011110000111011101110111011101110111100001111000011101110111011101111000011110010111100101111000011110000111100001111000011110010111101101111101100000011000110010010111100011101001100101111100100010010110101000101110001001010011000101101100011100010101000000111010010101110110111001101110010001110101000001110000011100110111001001110010011100010111000001101111,
	960'b011011000110110001101110011001100011100001001111011011100110111101101111011011110111000001110000011100000111000001110000011100010110101000101000001011110110000010001101100011001001011110010000100101101000011001111111011111110111101101111011011110010111100001111000011110000111100001110111011110000111011101110110011101110111100001111000011110000111011001110110011101110111011101110110011101110111011001110111011101010111010101110101011101100111010001110110011101100111011001110101011101010111011001110101011101100111010101110110011101100111010101110111011101110111010101111000011101110111100101111000011110000111011101110110011110000111011101110111011110000111100001111000011101110111011101111000011110010111100001111000011110100111101101111010011111101000001110010011100100001001011010001110011110011000000100111101001000110010011001101011011011100100110001000111011000100111000101110001010010100100100101110001011100110111001001110010011100100111000101110001,
	960'b011010110110110001101101010111010011001101011101011011100110111001101111011011110111000001110000011011110110110101110000011100010110010000101010010000100111101010001010100100111000101110000101100001100111110101111100011110110111101001111001011110000111011101111000011110000111100001110110011101100111100001111000011101110111100001110111011110000111100001111000011101100111011001110101011101100111010101110110011101100111011001110101011101010111011001110110011101010111011001110110011101010111010101110110011101100111011001110110011101100111010101110110011101010111011001110101011101010111011001110110011101100111011101110111011110000111011101110111011101110111011001110111011110000111100001111000011101110111100101111000011110100111101101111010011110100111101010000000100100001000101110010001100010011001011001011011001010000010011001101011011011110101011101011000011011010111010001110010010100100100010001110000011100110111001001110011011100100111000101110000,
	960'b011010100110110001101100010011100011010101100101011011100110111001101110011011110111000001101111011011010110110001110001011010100010111100101001010100011000001010000100100011101000011110000011011111100111101101111010011110010111101001111001011110010111100101111000011110000111100001110111011110000111011101111000011101110111011101111000011110000111100001110110011101100111011001110101011101100111010101110101011101100111010101110110011101100111010101110110011101100111010101110101011101010111011001110101011101100111011001110110011101100111011001110110011101010111010101110111011101110111011001110110011101100111011101110111011101110111011101110110011101110111011101110111011101110111011101111000011110010111100101111001011110010111100001110111011110110111101001111100100010001000010110001011100100011001100001101100001011110010100001101101011100010110010001101010011100010111010001110100010110010011111001101111011101000111001101110011011100100111000101110001,
	960'b011010010110110001101010001111100100000001101001011011000110110001101101011011110110111101101111011011000110111001110000011001110010000000101111011000101000100010000111100010001000001010001010011111000111101001111001011110100111100101111000011110010111100001111000011110000111100001111000011101110111011101110111011101110111011101111000011110000111100001110111011101100111011101110111011101100111010101110101011101100111010101110101011101100111011001110111011101010111011001110110011101100111011101110110011101100111011001110110011101010111011001110101011101010111011001110101011101100111011001110110011101010111100001110111011110000111011101110111011101100111100001111000011101110111100001111001011110000111100001110110011110000111100001111001011110000111101001111011100000001000000110001000100100111001000001110111001111000010110001101101011100110110110101110010011101000111010001110100010111100011100001101100011101010111001101110011011100110111001101110010,
	960'b011010010110101101100011001100010101000001101010011010110110101101101011011011000110110101101110011010110110111101110000011001110001111100110101011010011000101010001101100001111000000110001101011111010111101001111010011110100111100001111001011110000111011101111000011110000111011101111000011101110111011101110111011101100111011001110110011101110111011101110110011101100111100001111000011101100111011001110101011101010111010101110110011101100111011001111000011101100111010101110111011101010111011001110101011101010111010101110101011101010111011101110101011101100111011001110101011101100111011001110101011101100111011101110111011110010111100001110111011101110111100001111000011110000111100101111001011110000111100101111001011110000111101001111001011110100111100101111010011111101000000110001000100100111000110101111010010000100010111001101100011100110111001101110011011101000111010001110101011000100011010001101000011101100111010001110100011101000111001101110011,
	960'b011010010110101001010101001011100101110101101011011010010110100101101001011010010110101001101011011010100110111001101111011001100010000100111001011010111000101110010101100010011000010010001111011111000111110001111010011110110111100001111000011110000111100001111000011101110111100001110111011101110111100101111001011101100111011101110111011101110111011101110101011101010111011001110101011110000111011101110110011101100111011001110110011110000111011001110110011101100111010101110110011101010111011001110110011101010111011001110110011101010111011001110110011101010111011001110101011101110111010101110100011101110111011101111001011110000111100001111000011101110111011101111000011110000111100001111000011110000111100001111000011110000111100101111001011110110111101101111011011111011000010010001000100100101000110001111000010001110011000101101100011100110111001101110011011100110111001101110101011001110011001001100011011101100111010101110100011101000111010001110011,
	960'b011010010110011101000001001101100110011101101101011010010110100001101000011010000110100001101000011010010110100001011111010011110010001000111111011010111001000010100001100011111000100110010011100000010111110101111100011110110111100001111001011110000111100001111000011110010111011101111000011101110111100001111000011101100111011101110110011101110111011101110111011101100111010101110110011101010111010101110110011101010111010101110101011101010111011001110110011101100111011001110110011101010111010101110110011101100111011001110110011101010111011001110110011101100111011001110101011101100111011001110101011101110111100001110111011101110111011101110111011101110111100001111000011110000111011001111000011110010111100001111000011110000111100001111010011110110111101101111110100000001000100110001110100110001001000101110101010010010011011101101100011100110111001101110011011100110111001101110100011010010011010001011100011101100111010101110100011101000111010001110011,
	960'b011011110110011100110010010001010110110001101101011010100110100101101010011010010110100101100110011001100101110101011000010100100010001101000001011010011000111010100110100101011000110110010100100000111000000001111101011110110111100101111001011110000111100001110111011110010111100001111000011101110111011101111000011101110111100001111000011101110111011001110111011101110111011101110111011101000111010101110101011101110111011001110101011101010111100001110111011101010111011001110110011101110111011001110111011101110111011001110110011101010111010101110111011101110111011001110110011101110111011001110111011101110111100101111001011101110111011101110111011110000111011001111000011101110111011101111000011110000111100101111000011101110111100101111001011111010111111010000000100001001000110010010011100111011000111101110001010010100011101001101101011100110111001001110010011100100111001001110011011010110011011101010011011101000111010101110101011101000111010001110011,
	960'b011100010101111000101010010101100110111001101110011010110110100101101010011010100110101001100101011001000101111101100100010111110010011101001001011000011000010110101011101000001001010110010111100001101000001110000000011111100111101101111001011110010111100001111000011101110111100001111000011101110111100001110111011101110111011101111000011101110111011101111000011101110111011101110111011110000111011101110111011110000111100001110111011110000111011101110111011101110111100001110111011101110111011101110111011101110111011101111000011101110111100001110111011101110111100001110111011101110111100001111000011101110111011101111000011101110111011101110111011101110111100001110111011110000111100001111001011110000111100001111000011110010111101001111011011111111000001010000100100011001001001110011101101001111000011001101000010100100100001001101100011100110111001001110010011100100111001001110010011011010011110001001001011100110111010101110100011101000111010001110011,
	960'b011100000100110100101100011000110110111101101110011010110110100001101011011010100110100101100100011001100110011001100111011000010010110001010001010111100111110110100111101001111001110010010111100010101000011010000010011111110111101001111001011110010111100001111000011110000111011101111000011101110111100001110111011110000111100001110111011110000111100001111000011101110111100001111000011101110111100001111000011110000111100001111000011110000111100001111001011110000111100001111000011110010111100001111001011110000111011101111000011110010111100001111000011110000111100001110111011101100111100001111000011101100111011101111000011110000111011001110111011110000111100001111000011110000111100001111001011110000111100001111001011110110111101101111011100000001000010010000110100100111001100010100101101011111000000001100010010110000100100001101100011100100111000101110001011100010111000101110010011011110100010000111111011100000111010001110011011100110111001101110010,
	960'b011010110011011100110111011011000110111101101110011011000110100001101011011010110110011101100100011001110110011101101001011000110011001001011011011001000111010110011010101011011010001010011001100011111000100010000100100000010111101101111010011110010111100001111000011110000111100001111000011101110111100001111000011101110111100001111000011110000111100001111000011110000111100101111000011110000111100001111000011110010111100101111001011110010111101001111001011110010111100001111000011110100111100101111001011110010111100101111000011110000111100101111001011110000111100001110111011110000111100001111000011110000111011101110111011110000111011101110111011110000111100001111000011110000111100001111000011110000111100001111000011110010111101101111100100000001000010010001010100110111001111010101100101101100111100001100001011000110101000001101100011100010111000101110001011100010111000101110010011100000100110100110101011011000111010001110010011100100111001101110010,
	960'b010111100010100001001010011011110110111101101110011011000110011001101010011010100110001101100100011001110110011101101001010111100011100101101000011111100110100010000010101110001010110010100000101000001000110110000111100000100111110101111011011110100111100101111000011110000111100001111000011110000111100001110111011110000111011101110111011110000111100101111000011110000111100101111000011110010111101001111010011110100111101101111010011110110111101101111100011110110111110001111100011110110111101101111011011111000111101001111010011110100111101001111010011110010111100001111001011110000111100001111001011101110111100001111000011110000111011101110111011110000111100001111000011110000111100001111000011110000111100001111000011110110111101101111101100000111000011110010110101000001010100010111001101100100110110101110101011100010101101101101110011100000111000001110000011100000111000001110001011100010101011000101110011001100111001101110010011100100111001001110010,
	960'b010001010010011101101001011110110111101001111010011110000111001001110110011101100110111001110010011101000111010001110110011010000011110101100111100001100111000101110110101110011011001110100101101000001001010010001001100000110111110101111011011110100111100101111000011110000111011101111000011110000111100101111000011110000111011101111000011110000111100001111001011110010111100101111001011110110111101101111011011110110111110001111100011111010111110101111101011111010111110101111101011111010111110101111101011111010111110001111011011110110111101101111010011110010111100001111000011110000111100001111000011110000111100001111000011101100111100001111000011110000111011101111000011110000111100001111000011110000111100101111001011110110111101101111101100001001000110010011100100110111010111010111100100111110110101110000011011101000110000001101111011100010111000101110001011100010111000001110000011100010101111000101101010111100111001001110001011100010111000101110000,
	960'b001001010011111111001101110111101101110111011101110111011101110011011101110111011101110011011100110111001101110011011110110011100101101101011011011110011000101001101111100110101011101010101101100101101001100010010011100001000111110001111011011110100111101001111001011110010111101001111010011110100111101001111000011110100111101001111010011110010111101001111010011110110111110001111100011111010111111001111111011111110111111110000001100000011000000110000001100000111000001010000010100000101000000110000000100000010111111001111111011111110111111101111101011111010111101101111011011110100111100101111001011110010111100101111001011110000111101001111001011110010111100101111001011110010111100101111001011110010111100101111001011110100111101101111110100010111001100010010010100110101011011010100100011111101000010110000011011011000101110001110000011100100111001001110010011100100111001001110010011100100110010100101111010100110111000101110001011011110110111101101111,
	960'b000110010101100011011100111110101111100011111010111110101111101011111010111110101111101011111010111110011111100011111010110111010110111101011000011001100111110001111001100000111010111010110001100101111000111110010110100011100111111001111011011110110111101101111010011110100111110001111011011110100111101001111001011110110111101001111011011111000111101101111100011111000111110101111110100000001000000110000001100000011000000110000100100000111000010010000100100001001000010110000101100001001000010010000100100001001000001010000000100000001000000110000000100000000111110101111100011111000111101101111011011110110111100101111001011110100111101001111010011110100111101001111011011110100111101001111010011110110111101001111001011110110111110001111111100101001001000110010001100111101011000010001000011011111000101101110101011001000100110101101110011101000111001101110011011100110111001101110011011100110110101000110100010001110110111101110000011011110110111101101110,
	960'b000111110101000111011010111110011110011111011000110101111101011111010111110110001101101111011100110111101110011111111000110111100111100001001000010100010110001001110010011100011000111110101100100110101000111010001100100100111000000101111110011110110111101101111100011111000111110101111101011111010111110001111011011111000111110101111100011111000111110101111111011111101000000010000001100000101000010010000100100001011000010110000110100001111000011010001000100001111000100110001000100001101000011110000111100001101000010110000100100001001000001110000010100000001000000001111111011111010111111001111110011110110111101001111010011111010111101101111011011111010111110001111101011111100111110101111011011110100111110001111010011111000111111010000001100011001000101010010011100111111001011001110101011000000111011101100010010110010110110001110010011100100111001001110010011100100111000101110001011100100110110100111110001111100110110001110000011011110110111101101111,
	960'b001000000011011011010111111110111101100001000101001101110011101100111011010000010110000001101000011110111101110111111001110111110111100000100110001110010011111101000100010100100110011110000001101000011001101010001101100010001001000010001110100001001000000110000010100000001000001010000010100000101000000110000001100000000111111001111110011111111000000010000001100000101000010010000101100001101000011110001001100010001000101010001011100011001000110010001110100011011000111010001101100011001000110110001100100011001000101010001001100010011000100010000110100001011000010110000011100000100111111101111110011111100111111001111110011111111000000010000000100000011000001010000010100000011000000101111111011111110111110101111111100001111001000010001000100010101001001110011111100111110111000101011001011001000100110101000101001011010110110001110011011100010111000101110000011011110110111001101101011011100110110001001001001101110110100101110000011011110110111101110000,
	960'b000111010011000111010111111110111101011100110110001001100010101000101010001011000011001000101111010001011101100011111010110111011000000101101001001001100011010000110011010000000100100101101011100110101001110110010101100011101000100010010000100101001000111010000111100001101000011110001000100010001000011110000111100001011000010010000101100001011000010110000101100001111000100110001001100010111000101110001101100011101000111110010000100100001001000010010011100100111001001110010010100100101001001110010001100100011001000010001110100011111000110110001010100010101000100110000111100001011000010010000100100000111000001110000100100000111000010110000110100001101000100010001000100001111000011110000101100001001000001110010000100100001000011110000101100100101001110010011111100001010101010001010010010011100011111000110100011001010111001001110001011100010111000001110000011100000111000001101111011011110111000001010111001100010110001001110001011100000111000001110001,
	960'b000111010011000011010111111110111101011100110011001001100010101100101011001010010010100000100111001110001101011111111010110111011000001101110111001110110001010000100111001010100010110100111010011011101000001110011001101000011001100010010011100100111001000110011001100111111010000010011101100111001001110010011010100110001001100010010110100101111001011110011000100110011001101010011100100111011001111010100000101000001010001010100010101000101010001110100011101001001010010010100100101001001010001110100011101000111010001010100001101000001010000010011110100111011001110010011001100110001001011110010110100101101001010110010101100101101001100110011100100110111001111010011101100111001001110110011100100101101000111110001100100011101001000010011000100111111000110001110110010101110100001000111010001100100001110000100110011011100111010001110010011100100111001001110001011100010111000101110001011100010111001001100010001100010101100001110001011100010111000101110001,
	960'b000111010010111111010110111111001101011100110000001000000010010000100011001000000010000000100001001101011101011111111010110111101000010001111011011100100010010000010110001000000010011100101010010001000110011101111010100100011010000010011111100111111001111110011111101000001010000010011111100111101001111010011011100110011001011010010110100101101001011010010111100101111001101110011100100110111001110110100000100111111010000110100010101000101010010010100100101001001010010010100101101001001010010010100100101000111010001010100011101000001001111110011111100111011001101110011000100101101001011110010101100100111001010010010011100101011001101010011100100111011001111110100000100111111010000010011011100110011001100010011001100110101001101010011101100001100110110101010000001111110011100000110001001010110001110001100110011101010111010001110100011101000111001101110011011100110111001101110010011100100111001101101010001100110100101001110001011100100111000101110001,
	960'b000111100010111111010110111111001101011100110000001000000010001000011111000111010001110100011100001011111101011011111011110110110110001101010011011011110111000100110110000110100010001100100000001010000010111100111011010101000111110010010001101001111011011010111100101111011011101110111000101101111011010110110010101011101010101110101010101010001010011110101001101010101010110110101110101100001011000010110011101101001011001110110100101101011011010010110110101101101011011010110111101101111011011110110110101101101011010010110100101101001011001110110001101100001010111010101100101010011010100010100110101001111010011110101000101010111011000010110011101101001011011110110111101110001011011110110110101101111011010110110000100111111000011001110000010011110100001000110111001100110011000000100111001000000110011101110111011101100111011001110110011101100111010101110110011101100111011001110101011101010111011001110000001110110011111001101111011100110111001001110010,
	960'b000111110011000111010111111111001101011000101111000111100010001000100010000111110001111000011100001011111101011011111011110101110011100000100110001110100101011101010010000101100001100100100100001000100010010000101001001101110101011101101011011111001000111110110001110000011100011011001000110010001100011011000100110000011100000010111101101111001011111010111111101111101100001011000010110001001100010111000110110001101100011111001000110010011100100011001000110010001100100011001001110010001100100011001000110010001100011111000111110001111100011011000101110001001100001111000000101111111011110110111100101111001011110010111101110000001100001111000110110001101100101011001010110010101100100011000001101110101010110010000110011100010110000001010010001111100011001000101111001011010010010100011000011010000111100101111000011110000111100001111000011110000111100001111000011101110111011101111000011101110111100001110100010010100011010001101011011101000111001101110011,
	960'b000111100011000111010111111111001101011000101100000110100001111000011111001000000010000000011101001011101101011111111011110101110011001100100001001001000010110100110111001101000001010000011000001000000010000100100101001010110011110101000111010100010110000101111000100001011001000010011100100111111001111110100001101000111010010110100111101010101010110110101110101011111011001010110100101101101011100010111001101110101011101010111100101111011011110110111100101111001011101110111100101110111011101110111011101110111011101010111010101110011011100010110110101101101011010110110011101100101011000010101110101011011010110010101010101010101010100010100111101001011010010010100010101000001001101110001011011111100111000001011001010100110101001001000101001100110010110000101000001011100001100100011101011101000111110001111011011110110111101101111011011110110111101101111011011110100111101001111001011110010111100101111000010110010010111101100100011101100111010101110101,
	960'b000111010010111011010110111111001101011100111100001011000010111100101111001100000011000000101111001111101101011111111011110101110011001100100010001001100010101000101111001110000011001100011101000100010001111000101011001010010010100000101001001011000011001000111110010010000100110101001111010011100100111001001111010011010100110001001100010010010100100101001001010010100100100001001010010010100100110101010010010101010101101001011101010111110110000101100000011000100110001001100101011001000110010001100100011001000110001001011101010110110101100001010110010101000101000001001100010010100100100101000110010001000100010001000011010000110100010101001001010010110100110101001101010011010100110101001100010010100100000000110000001011100010111000101011001100000010100100010011000111110110110101110110011111010111111001111110011111010111110101111101011111010111110101111101011111000111110001111011011110110111101101111011011001010010110101011000011101110111011101110110,
	960'b001000110011000111010111111110101110011111011000110101101101011011010110110101101101011011010110110110001110011111111010110101110011000100100011001010100010101100101100001101010011011000110101000100110001000100010110001001000010101100100111001001100010101100101111001100010011001100110101001101010011010000110011001100000010110100101011001010100010101000101010001010100010101100101100001010110010111000101111001100010011010000111000001110000011101000111100001111100011111000111111001111010011110100111100001110100011100100110111001101100011010100110001001011110010110100101110001011000010101000101010001010100010101100101011001010110010110000101110001100000011001000110011001100100011010000110010001100110011000000100111001001000010101000101111000111000001100000011110011100011000001110000010100000011000000110000001100000001000000010000000100000000111111101111111011111100111110101111101011111010111110101111101011011110011000001001001011101110111100101111000,
	960'b000111100010111111011000111111001111100111111011111111001111101111111011111110111111101111111011111110111111100111111100110110000011001100100010001010010010100100101000001011100011010000110111001110000011001100100000000101100001000000010110001001010011110101001111010010110100011001000100010001010100010001000100010000010100000101000010010000100100000101000000001111100011111101000000001111110100000101000011010001000100010101000111010010100100101101001110010100000101000101010001010011100100111101001110010011000100101001001000010010000100010001000101010001010100010001000011010000010100001001000001010000100100001101000100010001110100100001000110010010000100110101001101010010110100101001001100010100110101100000111110000111110001000100001110001000110111010001111101100001011000010010000100100001011000010010000100100000111000001110000011100000101000001010000010100000011000000110000000100000000111111110000000011101110011100000111011011101100111101101111001,
	960'b000111010010111011000110110110011101011111010111110101111101011111010111110101111101011111010111110101111101011111011001110001110011001100100100001001100010010100101001001011010011001000110100001101100011100000111000001110110001100000010000000011110001010000101101001111010100010101010011010010110100010101000111010100000100111101000100010000010011111100111111001111110100001100111100001111010011111001000000010000100100010101001111010010100100110001001111010100010101001101010100010110100101000101001111010011010100100101000111010001100100101101000100010000100100000100111111001111100100000001000110010000010100000001000001010000100100010001001110010011110100011101000110010011000101000101000100001111110010111100010011000101010000111100100000011101111000101010001001100001111000011110000111100010001000011110000110100001011000010110000110100010001000010010000100100001001000010010000011100000111000001010000010011111100100011000110001011100100111110101111011,
	960'b001000100010001000101111001100100011001100110100001101000011001100110011001100110011001100110110001100110011010000111010001101110010100000101000001001010010011000101011001011010011011100111000001100010011001100111001001111000011111100101000000110000001001100010010000100100001111110001010010011010001001100011101011110110111001100011111000101100001011100011000001101010101010100011101000110010001101000011010000110010010111101100010001000000001101000011011000111000001101100101011011011100010011000011011000110110001110100011011001001110110111000101010000110100001101100011011000110100010011001101110001010110001101000011011000110110010101010000010011110010010000100010110010111001001000000100101000110010001100000100010011100100100100001111101100011001000101110001011100010111000101010001010100010111000101010000110100001101000100010001000100010001000011110001000100001111000011110000110100001101000010110000110100001010101100100101110011011001000000001111110,
	960'b001010000010000100011111001000010010001000100100001001000010010000100101001001000010010000101000001001110010011100101010001010100010100100101010001001000010100000101001001010110011011100111100001101000011011100111110001110000011010100110111001110110011101000111000001110000011111001001001001111110011011000110110001111100100010001000001010011010101111001100011011000110110110001101000011001100110101001100111011000010110010101101100011001100110011001101001011010110110110001101111011101110111001101110011011101110111100001110111011110011000000001110101011101000111010001110110011101010111100010000000011110010111010001110100011101110111100110000101100010100111110100111100010110001001010010001100100011001000110010010000100111011001101010011111100111101001111110011111101000001010000010100001101000011010000110100000101000001010000110100001101000001001111110011110100111011001110010011011100110101001100110011001100110000111000000101011011011001001001110010010,
	960'b001010100010011000101000001010010010100100101001001010100010110000101101001011010010111100110100001101010011000100110010001101100011010000110100001011010010110000101011001100000011011100111010001101110011100100111111001111100011110000111110001111110100000001000001010000100100010101000111010011100101000101001101010011000101011101100010011100110111111110000000011111000111101001111010011110001000000010000011100000101000010010000100100001011000100110001100100011111000111110010001100100111001100010011011101011011010111110100010101000011001111010100001101000101010001110100100101001001010011010100111101010101010100110101010101011111010111110101110101101101011010001011001010111011011011111000000101111011011110010111100101111001011110110111100101111001011110110111101101111011011110010111100101111001011110010111100101110111011101010111001101110001011010110110010101100001010111110101101101011001010101010101000101001111000011000101110011001011010001110100100,
	960'b001100000011001000110100001100100011001000110100001101010011010100110101001101010011011000110111001110000011100000111010001110110011110000111100001110010011101000111110001111110011111001000001010000010100001001000111010010110100101101001100010100010101010001010110010111000110011101101100011100010111010001110100011101010111011001111000100000001000001110000000011111100111110001111011011111101000001110000101100001101000011110000110100001111000100010001010100011011000111010011000101000111010111010110001110101101101111111000011101111011011111011000000101111101011110010110111101111001011111110111111110000011100000011000000101111011011110110111010101111011011101001100110010100101011100010111110101110111011101010111010101110111011101110111010101110111011110010111100101111001011101110111011101110111011101110111011101110111011101010111001101110001011011110110110101101011011010010110011101100111011001010110000101100001001100000110110010101011010100010101110,
	960'b001110010011110000111111010000100100001101000100010001100100001101000011010001000100001101000010010000010100000101000011010001000100010001000110010001100100100001010000010101100101010101010010010100100101010101011001010111010110010101101011011101000111100101110111011110000111110110000011100000111000010110000101100001111000100010001001100011001000111110001100100010111000101110001101100100011000111110010010100101111000111110001101100101001000111010010010100101001001100110100100101011001011000110110111110111011110100011001001110000111100010011000010110000101100001111000011110001011100010011000100110001001100010011000011101101101011011010111000101101111011010101110100010001001010111010110110101100111011000110110000101100011011000110101111101011101010110010101010101010101010100110101010101010011010011110101011101011001010101110101001101001111010011010100110101001101010011110101000101010011010101010101011101011011001110100111111010010101010100110110100,
	960'b010011000100110101010001010101010101100001011011011000000110000101100001011000100110001001100001011000000110001001100100011001000110001101100100011001000110010001100110011010010110101001101010011010110110111001110001011101010111101101111110100001001000010110000101100001011000011010000110100010001000100110001001100010111000110110010000100101001001010010010001100011011000100110000101100000010111010001111001100010011000111010100100101011101010110010101111101100001010111010101111101100001011001010111000110110011110001011000100101111111011101110100101101001111010111010111100110000111100000111000000110000001100000011000001110000001100000011000001110000101100001110001011001111011010100111000000101111001011101110111010101110011011100110110111101011011000111010001100100101111001010110001011100010011001010110010101100100111001110010011000100101011001010110011101100111111001111110011111100111011001101010011100100111001001010001001001001110011001010110100011,
	960'b011010010110100001101001011011000110111001101110011100010111010101110111011110010111101001111011011110110111110001111101011111010111110101111101011110110111101001111010011110100111101001111100100000001000000110000010100001001000011010000111100010011000100110001001100010101000101010001001100010001000100010000111100010011000110110001101100011011000100001111110011101110111010101110000011100010111001001111100100011001001100010100010101001011010001110100010101001001010001110100011101000111010101110110100101110111011111110110011101100011011010010110001101100111011011010111100101111111011110010111010101110001011100010111001101110011011100110111001101110011011100010001110001110001001101110111000101101001011010010110100101100101010110110100110100101100111100001101101011011100110101101100110011001010110011101100110011001110110110001101000011001110110011101110011011110100111100001110101011011110111000001111000011111000111111001001010001011010111111010010010,
	960'b100001001000010010000100100001011000010110000011100000111000010110000101100001011000010010000100100000111000001110000100100000111000001010000010100000101000001110000011100001001000010010000101100001101000011110001000100010011000101010001011100010111000110010001110100011101000111110001100100010001000100010001000100001111000011001111011011101000111000101110010011100110111010001110011011101000111010101111000011111101000101110010100100111001001110010010000100010101000110010001010100001111000110010010001100100001001000010001111100011101001011010011001100110101001111110100001101001101010100010101010101001111010100110101011101010101010011110100101101000111010001010000111001100111000001110100101101000011010000010100010100111101001101110011010100101001000100110000101100001101000001110000011011111000111011001110001011011000110100001100100011000100110001001100001011000100110001001100001011000110110001001100000011000000101111001000010001001000101101001101110,
	960'b100000001000001010000101100010011000100110001010100010111000110010001101100011001000100110000111100001101000011010000111100001101000011010000111100001111000011110000111100010001000100110001000100010001000100010000111100001111000110010001110100011101000110110001000011111110111101101111010011110100111110001111000011101100111101001111000011101000110111101110101011110010111101001111000011110000111100101111010011111011000000010000001100001011000100010000100100000111000101010010011100011101000011110000111100100101000110110000111100010001000011110000001100000011000010110000101100010001000101010001101100100001001010010010110100110001001100110011001100110011001100110000110001101010110110110010001100011001000110010001011100011011000111110010000100011011000101010001010100011101000110010001110100100011001000110001001011111000111101101111000011110110111111101111111100000011000000010000000100000011000010010000110011111100111010101010011001000110101110001111010,
	960'b100000011000000110000010100000111000010010000101100001101000100010000010011101110111001101110010011011110110110101110011011101100111011101110111011101110111011001110111011111011000001110000001011110010110111101101101011111011001001010010110100100111001000110001100100000010111010101110010011110011000001001111100011111010111101101111100011101110111000101111011100000111000010010000001100000101000010010000100100000111000001110000110100001101000100010001011100010111000110110010101100101111001001110010101101011001010011110010110100101001001001010001100100000111000000001111110011111110111111110000000100000101000010110000100100001101000011110001010100010111000100101111001001101010101010101111101011110110111101101111011011110100111101101111110011111010111101001110111011101110111100101111001011110100111101101111001011101010111010001110011011101010111100001111010011110110111110001111110011111111000010010000101100000000111110001011111001000110101010001111011,
	960'b100000011000001010000011100001001000010110000101100001011000010001111011011010000101100101001111010010100100011101001001010011000100111101010101010110000101011001011100011011010111100001110111011011100110001101100110100001001001010110011000100101111001010110010000100000100110011101100100011011000111100101111000100000111000001110000010011111000111011110000001100010101000101110001010100011001000111110001101100011101001001110010111100101011001100110011100100110011001100010011100100111111010000110100111110011001100100110101011101001111010010110100001100110101001001110001101100001101000010010000001011111100111011101110100011101010111010101110111011110000111011101101111001110000100100001110100011101000111000101110001011011110110111101110000011011110110110001101011011010100110111001110000011100100111000101101111011011100110111001101111011011100110111101110011011101100111011001110111011110000111011001110101011101000111010001011110001000110100100001110110,
	960'b011111101000000010000010100001001000010010000101100001011000010110000110100001000111111101110010011000110100111101000110010001100100100001001111010100110101011101100000011011100111011101111101011110100111011101111100100001001000001010000010100001101000101110001100100010000111011001110001011110101000110110001011100100011001000110001111100001100111111110001001100100011001001010010001100100011001000110010010100101001001011010010111100101111001011110010101100101111001101110100000101001011010100110110000110101101101010010110000101001101010000110011110100111011001110010011100100110111001100010001111100001010111110001111001011100110110111101101111011011010110101101100110001110000011111001101011011010110110011001100101011001000110001001100001010111110101111001011111010111110110000001100011011001010110011101100111011001110110011001100111011010000110101101101110011100000111001001110100011101000111001101110000011011110110111101011100001001000100001001110010,
	960'b011110110111110001111100011111010111111001111111100000001000000010000001100000101000000101111010011100010110100001100000010110100101010001010100010101100101111001101100011100000111010101111000011101100111000001101011011011100111101010000110100010101000110110010000100100011000110110001010100100001001110010011011100101011001011010011011100110001001001010010101100110111001101110011000100101101001011010010111100101111001100010011000100101111001011110010110100110111010000110100101101010101010110010110010110101011101011010110111101011101010101010101000101001111010100110101100101010001010001110011111100111011001011010001101100001101000000101111111011110100111011001101111010000010011100001101011011010010110000101100000011000000101110001011001010101110101010001010011010101010101011101010110010101100101100101011011010110100101100001011010010111000110000001100000011000110110011101101010011010110110101001101001011010000110100001010111001000010011110001101010,
	960'b011111100111110101111100011110110111101001111011011111000111101101111010011110100111101001111011011111000111110001111100011111000111101001111000011101100111001101101110011001100110001101100000011000000110000001011101011000100110111101110111011111000111111110000000100000101000001110000010100001001000011110001001100010101000110010001110100100011001000010010110100110001001100010010100100110101001101010011001100111001001111010100000101000111010000010011101100111111010001110100110101010101011000010111001110110011101101010111011101100101010111010101110101011011010110010101011101010011010011110101000101011101010110110100100100111011010000010011111100110011001001110001011010101100011011101111001011111000111100001110011011010110110011101100001010110110101011001010100010101010101011001010101010101000101001101010100010101000100111001001100010011010101000001010011010101110101101001011011010111010101110101011101010111100101111101010000001000010011100001100001,
	960'b011111000111110101111101011111010111110101111101011111010111110101111101011111000111110001111100011111010111110001111100011111010111111001111101011111100111111101111111011111100111101101111000011101010111000001101001011000100110000101100001011000010110010101101100011101010111101101111110100001001000100110001111100101111001011110010010100011001000011110000001100000001000001110001010100011011000100110001010100011111001010110011001100111111010000010100011101001011010010110100101101011001011010110111111110111001101101010111010101101001011000110101111101011011010110010101101101011101010111010101101101011011010011110100100100111111001111110100100101001001010001010100001011011100011100010010000101000011001110010010101100011101000110110000110011111000111011101110010011100000110111101101100011010010110011101100111011000110101110101011000010101010101001101010011010100010100111101001110010011100101000101010001010101010101011101001000001000000011010001011011,
	960'b011110110111101101111011011111000111110001111101011111010111111001111101011111100111111001111111100000001000000010000000100000001000000001111111100000001000000110000010100000101000001010000010100000101000010010000100100001001000000101111101011100100110010101100010011001010110011101101101011100010111100010000001100100101001111110100110101001111010011110100001100110011001010010011000100110001000101110000100100001001000010010000101100010101000110110010010100110001001011110011000101000011010100010110010110011111100110110111000101101101011001110101110101011011010101110101010101011001010110110101101101011111010111010101101101011001010110110101101101010101010011110100110011111000011100010010010101001001001110110011011100110111001111010011011100101001001001110010100100011111000011010000010100000001000000001111001011011100110101001101110011011110110110001101001011001000101111101011100010101110101001101010000010100000101000001000011001000000011000001010100,
	960'b011101100111100001111001011110100111101101111100011110110111110001111101011111100111111001111111100000001000000110000001100000011000000110000010100000101000001110000100100001001000010010000101100001001000010110000101100001101000011010000111100001111000010110000010011111100111100001110110011100000111000101110001011100000111011010000010100010011001010110100011101010011010001110100001101000101001110010011001100101111001010010001111100010011000100010000101100001011000010010000101100010101001001010011000101000101010101010101010101010011010100010101001101011011010101110100101101001101010100110101011101011001010110110110000101100101011001010101111101011011010110010101110100011000011100010010000101010101010010110100100101001101010011110100011100111111001110110011010100110011001010010010000100011001000100110000111100000100111111101111111100000000111110101111010011110000111100001110110011100010110110001100110011000100110000101010010001000100011001001011110,
	960'b011010110111001001110100011100100111001001110100011100100111001101111001011110100111101001111010011111000111110101111101011111010111111001111110011111100111111110000001100000111000001110000100100000111000001110000100100001011000010110000110100001101000011010000110100001101000100010001000100010001000100010000111100000110111111101111101011111011000000110001110101010011010111110101011101100101011001010101111101010101010011010100011101000001001111010011000100011111000100110001000100001111000101010001011100010001000101010010001100101011001001110010100100101101001110110100101101000011001110010011111101000101001111110011111101000101010101010101101101010011010000110100110100011110011010110000010101010001010001110100000101000101010010010100011101000011001110110011001100110111010000010011011100110101001100110010111100101001001001010001110100010001000011110000101100000111000001110000100100001001000000110000000011111110111110001100111001001010011010101101110,
	960'b011001110110101101101010010111100101111101100110011010000110110101110010011100100110111101110000011101000111011001111000011110010111101001111011011110110111110001111101011111111000000110000010100000111000001110000100100001011000011010001000100010011000100110001001100010011000100010001001100010101000101010001011100011001000110010001010100010001000100110010011101001011010110010101111101101011011100110111010101110011011101010111000101110001011100010110111101101011011000110101010101000101001111110011101100101101001001010010011100101011001000110000111100000111000100010001101100011001000100110001010100010101000011010001000100011001001010110011010100111011001011110010111100001100011001101110100101001001010000010011100100111011010001010100011101000111010000110100100101001111010100110100100101000001001111110011001100101001001000010001111100011101001001110010010100011111001000110010000100011011000100110001000100001111000011101101110001001110011100101110011,
	960'b011011010110101101101010011010110110101101101100011010010110110001110001011100000110101001101010011100000111001101110100011101100111011001110111011101100111011001110111011110100111110001111101100000001000001110000101100001101000011110000110100001111000011110001000100010101000101010001011100010101000101010001011100010111000101110001100100011001000111110010100100110001001101110011111101000111010100010101101101100001011011010111000101101111011100010111000101110001011011110110101101100111011000110101111101011101010101110101001101010001010010010010011100010111000011110000011100000101000000001111101011110100111101101111111100001101001000010001001100010001000100110001011011111110011010001011111100011111000101110000101100010011001010010011100101000001010000110100001100111001001100110011001100100111001001110011001100110111001011110010110100101011001010010010001100100111001100110010111100101011001011110010110100100111001001001110100001001100011110101111000,
	960'b011011010110100001100110011010010110101101101110011011000110111001110011011101000111010101110110011101100111011101110110011101100111011101111000011101110111011001110101011101000111011001110111011110100111111010000001100000111000010010000001100000101000001110000110100010001000100110001001100010011000011110000111100010101001001010011001100111101010010010101001101011001010111010110001101101001011011010110110101101011011010110110110101101011011010010110100101100111011010010110100101100111011000110101101101011101010110010101100101011001010101110100111101001001010001010011111100101111000110110000011011111010111101101111000011110010111111001111100011111101000000110000011011110010011001101001111011111111000000110000000100001001000100010001010100011001000110010001101100100111001100110011001100100111001000110010100100101111001100110011010100111001001110110011001100110001001011010010110100101111001100010011000100110001001011101110101001000010011110001111111,
};
parameter [0:85][959:0] b_picture = {
	960'b011100000111011001110111011110000111011101101111011000000101001001000101010011010110111101111000011110010111100101111010011110100111100101111010011110100111100101111010011110110111101101111011011110110111101101111011011110110111101101111010011110110111101001111010011101100111011001111001011111100111111101111111011111110111110101111001011110000111100101111001011110110111111010000000100000000111110101111111100000011000010110001000100001101000000110000010100001111000111110010011100011111000110110001011100010101000100110001000100001011000001010000001100000000111111101111110011111100111110101111100011111000111101101111011011110110111101101111010011110100111100101111001011110010111100101111001011110010111100101111001011110010111101001111010011110010111100101111001011110010111100101111001011110010111100001111000011110000111011101111000011110000111100001111000011101110111011101110110011101110111011001110110011101100111011001110110011101100111010001110100,
	960'b010001110101100001101111011100100111001001101100011000100101001101000100010010000110011101110010011100110111001101110100011101000111100001111001011110010111100101111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111100001110101011101000111011001110111011110000111101101111100011111000111110001111001011110100111101001111001011110110111111010000001100000111000001010000011100001101000100110000110100000110111111110000000100001101000101110001101100010101000100010000110100001001000001110000001100000001000001110000010100000000111111101111110011111010111110001111100011110110111101001111010011110100111100101111001011110010111100001111000011110000111100001111000011110000111100001111000011110000111100001111001011110000111100001111000011110000111100001111000011110000111100001110111011101110111011101110011011100100111001001110010011100100111000101110001011100010111000101110001011100010111000101110000011100000111010001110100,
	960'b010001010011111001000110010010000100100001001000010001110100011001000100010001000100011101001000010010000100100001000111010010110111010001111001011110010111100101111001011110010111101001111010011110100111101001111010011110010111100101111001011110000111010001110011011101010111011001110110011101110111101001111010011111000111110001111100011111000111110101111100011110110111101101111101011111101000001010000110100010001000010001001110010010010100100101001001010010100100101001001010010010100100101001001010010010100100101001001000010011010111111110000011100000010111111101111110011111010111110001111100011110110111101001111010011110100111100101111001011110000111100001111000011101110111100001110111011101110111100001111000011110000111100001111001011110000111100001111000011101110111100001111000011101110111011101110111011110000111001101001011010001110100100001001000010010000100100001001000010010000100100001001000010010000100100001000111010010110111000001110101,
	960'b010101010100101101000100010010110100110001001100010011000100110001001100010011000100110001001011010010110100110001001010010001110111001101111001011110000111100001111001011110010111100101111010011110100111100101111001011110010111100001111000011101110111011001110101011101010111011001111000011110000111101001111100011111000111110001111100011111010111111001111111011111010111110001111101011111101000000010000101100010011000001101001000010010100100101101001010010010100100101001001010010010100100101001001010010010100100101101001010010010000111111110000100100000011000000001111110011111010111110001111100011110110111101001111010011110010111100101111001011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001110111011110000111011101110111011101110111100001110111011101100111010101110110011101110111001001000111010010110100110001001011010010110100101101001011010010110100101101001011010010110100110001001011010001110111000001110101,
	960'b010111110101000001000101010011000100010101000011010001000100010001000011010000110100010001000110010010000100010101001011010010000111001001111000011110000111100001111000011110010111100101111001011110010111100101111001011110000111100001111000011110000111100001111000011110000111100001111001011110010111101001111010011110110111101101111010011110110111110001111101011111100111111110000000100000011000001010000101100010001000001101001010010010110100010101001001010010100100101001001100010010110100101001001010010010100100010101001011010010010111111110000100100000011000000001111110011111010111110001111011011110100111101001111001011110000111100001110111011101110111011101110111011101110111011101110111011101100111011101110110011101110111100001110111011101110111011101110111011101110111011101110101011101000111001101110101011101100111000101001000010011000100010101001000010010000100100001001000010010000100100001001000010010000100010101001100010010000111000001110101,
	960'b011001010101011101000110010011000100001100111000001111100100001100111001001100110011101101010110011001110100011101001011010001110110001001101101011010110110011001100101011010100110110101110100011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100101111001011110010111101001111001011110100111101101111100011111010111111001111111100000011000001110000011100001101000001001001010010010100100100110000001100011011001101010100110100111111001000110001100100000110100100101001010010010010111111110000100100000011000000001111110011111000111101101111010011110100111100101111000011110000111011101110111011101100111011001110110011101100111011001110110011101100111011001110110011101100111011101110111011101110111011101110110011101100111011001110101011101000111001101110011011101010111000101001000010010110100100001101101011100010110111101101110011011110110111101110000011010110100100001001011010010000110111101110100,
	960'b011010000101111001000110010011000100001100110011001101100011100000110011001011010011001101000011010011010100010101001100010001010100110001000100001111110100011101001100010100000101100001011101011011000111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001111001011110010111100101111001011110100111101101111100011111000111110101111110100000001000001010000010100001011000000101001010010010100100100110001011101100111101010011011011110101001011011010010010100001010100101001001010010010010111111110000011100000010111111101111110011111000111101101111010011110010111100001111000011101110111011101110110011101100111011001110110011101100111011001110110011101100111011101110111011101110111011101110111011101100111011001110110011101100111010101110101011101100111010101110100011101010111000001001000010010110100100001110000011101010111010001110011011101000111010001110101011100000100100001001011010010000110111001110010,
	960'b001111110100111001000110010011000100001000101010001100100011000000100111001001100010110000110000001101000100001101001101010000110011010000110001001110010100010101010001010101000110011001100110010110010110110101110110011101100111011001110111011101100111011101110111011101110111011101110111011110000111100001111000011110010111100101111001011110100111101001111011011111000111110101111110100000001000000010000010100001001000000001001001010010100100101010011011110110001110000011011101110111001101001010011101100000100100100101001010010010010111111010000011100000010111111101111101011111000111101101111010011110010111100001110111011101100111011101110110011101100111011001110110011101110111011101110111011101110111011101110111011101110111011001110110011101100111011001110101011101100111011001110101011101010111010001110011011100100110110001001000010010110100100001110000011101000111001101110010011100110111001101110100011011100100100001001011010010000110110101110001,
	960'b001001100010101101000010010011010100000100100101001010010010110000100000001000100010101000101101001011110100001001001101010000110011011000111101010000010101000101011110011000010110100001110100011011000110011001110011011101100111011001110110011101100111011001110110011101100111011101110110011101110111011101110111011110000111100101111000011110000111101001111010011111000111110101111110011111111000000010000001100000110111111101001001010010100100110010101010111000101110000111011101110111001101100110100111100000010100100101001010010010010111111010000010100000000111111001111101011111000111101101111010011110010111100001110111011101100111011001110110011101100111011101110110011101110111011001110111011101110111011001110101011101100111011001110110011101100111010101110101011101010111010101110100011101000111001101110010011100100110110101001000010010110100100001110000011101010111010001110011011100110111001101110011011011000100100001001011010010000110110001110001,
	960'b001001000010010101000001010011010100001000100111000111110010000100011111000111110010010000100110001010010100001001001101010000110011011101000010010010110101101001101010011100010111000101110101011101110111001101110100011101010111010101110101011101100111011001110110011101100111011001110110011101110111011101110111011101110111100001110111011110000111100101111010011110100111110001111100011111100111111110000000100000110111111101001001010010100100110010100110111001001110010111011111110111111101100110100011100000100100100101001010010010010111111010000010011111110111110101111100011110110111101001111001011110010111100001110111011101100111011001110110011101000111001101110101011101100111011001110110011101100111010001110100011101010111010101110101011101000111001101110101011101010111010101110100011101000111001101110011011101010111000001001000010010110100100001110001011101010111010001110011011100100111001001101011010111000100011001001011010010000110110001110001,
	960'b001111100011001001000010010011010100000100100001000111000001110000011100000111010001111100100010001010100100001001001101010000110011100101000101010101100110100001110010011101010111011001110111011101100111011001110110011101010111010101110110011101100111011001110110011101100111011001110110011101100111011001110110011101110111011101110110011101110111100001111001011110100111101101111100011111100111111110000001100000110111111101001001010010100100101010010010110100001110011011100100111000011100100110010100100000100100100101001010010010010111110110000001011111100111110101111100011110110111101001111001011110010111011101110101011101000111010101110011011100010111001001110011011100100111010001110101011101000111010001110101011101100111010101110101011100110111001101110011011100110111010101110100011101000111010001110100011101010111000101001000010010110100100001110001011101100111010001110010011100100110000101001101010100000100010101001011010010000110101101101111,
	960'b011000010100110001000101010011010100000100100000000111000001101100011011000111100001111100100011001010100100001001001101010001000100000001001100011000110111001001110110011101100111011001110110011101110111011001110110011101100111011001110101011101100111011001110101011101010111010101110110011101100111011001110110011101100111011101110110011101110111100001111001011110100111101001111011011111010111111001111111100000100111110001001001010010100100100110000110100111111100011111010111110001111001111110001011100000100100100101001011010010010111101101111111011111010111110001111011011110100111101001111001011101100111000101110001011100000111000101110001011100010111001001110011011100110111010001110101011101000111010101110101011101010111010101110100011100110111001101110011011100100111001101110100011101000111010001110101011101100111000101001000010010110100100001101111011101010111010001110011011011000100100101000100010100000100011001001011010001110110100101101101,
	960'b010010110100011101000101010011000100001000101001001000100001111100100100001000110010001000100101001010010100000101001101010000110011100001000110010111110110111001110101011101100111011101110111011101110111011001110110011101010111010101110101011101010111010101110101011101010111011001110110011101100111011001110110011101100111011001110110011101110111011101111000011110010111100101111010011110110111110001111101011111110111101001001001010010110100100101111100100001001000101010010000100010111000010010000011011110110100100001001011010010010111101001111110011111000111101101111010011110010111100101111001011100110111000101110001011100010111001001110010011100110111001101110100011101010111011001110110011101100111011001110101011101010111011001110101011101010111001101110010011100100111001001110010011101000111010101110101011101010111000001001000010010110100011101100000011011100111000001101101010111100100001101000101010011110100011001001011010001110110010101101010,
	960'b001001010010100001000001010011010100010101000010010000010100000101000001010000010100000101000001010000100100010101001100010000100011010000111100010001110100110101011011011010100111000001110100011101100111011001110101011101000111010001110100011101010111010001110011011100100111001001110100011101010111010101110101011101010111010101110101011101100111011101110111011110000111100001111001011110100111101101111100011111100111100101001001010010110100010101001001010010010100100101001001010010010100100101001010010010010100010101001011010010010111100101111101011110110111101101111000011100100111010001110101011100010111000101110001011100110111010001110011011100110111001101110100011101010111011001110110011101100111011001110101011101100111011101110111011101100111001001110010011100100111001001110011011101010111010101110101011101100111000001001000010011000100010101000110010010000100100001001000010001100100010001000100010001010100010101001100010001110110001101101010,
	960'b001010000010101001000010010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001100010000110011100101000001010011000100101101001100010110000110010001101010011100000111010101110011011100110111001101110011011101000111010001110001011011110110111101110010011101010111011001110110011101100111011001110110011101110111011101110111011110000111100101111001011110100111101101111011011111100111100101001000010010100100101101001011010010110100101001001010010010100100101101001011010010110100101101001010010010000111100001111100011110100111100101110110011100010111001001110011011100100111000101110010011100110111010001110100011100100111001001110011011100110111010001110110011101100111011001110110011101100111011101110111011101010111000101110010011101000111010101110101011101010111011001110110011101100111000001001000010010110100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010001110110001001100111,
	960'b010001010100011101000100010000100100001001000011010000100100000101000001010000010100000101000010010000100100001001000010010000100100000101000001010000100100001001000111010100110110000001101001011001100110111001110011011100110111001001110010011100110111010001110001011011100110111001110000011101010111010101110101011101010111011001110110011101110111011101110111011101110111100001111001011110010111101101111011011111010111100001001100010001110100100101001001010010010100100101001001010010010100100101001001010010010100100101001000010011000111011101111011011101110111001101110010011100100111001001110101011101000111001001110010011100100111010001110011011100110111001001110011011101000111010101110110011101100111011001110111011101100111011101110111011101100111010001110101011101100111011001110110011101010110111101100101010111110101100101000100010001000100011001000110010001000100001101000100010000110100001101000100010001000100010001000100010010010110010101100101,
	960'b010111110101101001000100001011000010011100101111001010110010000100011100000111000001110100100110001010100010101100110001001110000100001001001111010011100100010101000000010000110101000001101000011011010110110101110010011100100111000101110000011011110111000101110000011100000110111101101100011011010111001101110100011101000111010101110101011101100111011001110110011101100111011101111000011110010111100101111010011110110111101101111000011101110111011101111000011110010111100101111001011110010111100001111000011101110111011001110110011101100111100101110101011100100111001001110010011100100111010101110101011101010111010001110011011100110111010001110011011101000111001101110100011101010111010101110110011101100111011001110110011101110111011101110111011101110111011101110111011101110111011101110110011011110101111101010001010000110011101100111000001111100100101101001111010001000011100100111111001110010011011100111100001111110100001001001101011000000110010101101001,
	960'b001110110010110100100010000111110001111100100011000111100001100100011000000110000001101000100010001011010010111000110000001100110010111000110110010010000101010101011001010101100100101001011000011011100111000101110010011100100111001001110001011011110110110101101000011010100110111101100010011000100110111101101011011100100111011001110110011101100111011001110110011101100111011101110111011110000111100101111001011110100111101001111011011111000111110001111101011111100111110101111101011111010111110001111100011110110111101001111001011110000111010001110001011100010111000001110000011100010111001101110100011101000111010001110011011100110111000101101100011011000111000101110100011101000111001101110010011100110111010101110110011101110111011101110111011101110111011101110111011101110111011101110110011100110110111101101001011000010101010101000100001100100010110100110111001111100011010100110000001100000011000100110101001101110011111101010010010111010110001001100110,
	960'b001000000010001000100100001010110010110000101000001000000001101100011001000110010010000000100111001101000100100101001000010011000100000000110111001110100100101001011001011001100101111001001011011000000110111001101111011100000111000101110001011011010110011001100011010111110110011101011110010110110110001001101011011101000111010101110101011101100111010101110101011101100111011001110110011101100111011101111000011110010111101001111001011110100111101001111011011110110111101101111011011110100111101001111001011110000111011101110110011101000111010001110010011100010111000101110000011100000111000101110010011100100111001101110010011100100111000001100101010100010101100101101010011100000110011101011100011001010111001101110100011101010111011001110110011101100111011101111000011110000111100001110111011101110111011101110111011011110101110001001100010000000011000000100110001010000010100100100110001010000010110100110010001100110011111001001101010101000101011101010100,
	960'b001010100011000100111100010001100011001100100010000111110001110000011011000110110010101101000000001011110011110001000111010100000101110001001101001111010011111101010000011000010110101001011011010101000110001101101100011011100111000001101110011011000110101001100100010110100101010001010011010100010101100001100011011010100111001101110110011101010111010101110101011101000111010001110101011101010111001101110101011101100111100001111001011110000111100001111001011110100111101001111001011110000111100001111000011101110111011101110111011101100111010101110011011100100111001001110001011100000111000001110000011011110111000001110001011100100111000101100110010010110011111001001000010110100100101101001011011001010111001001101101011011100111001101110100011101000111010101110111011110000111100001111000011101110111100001110111011011100110010101011101010100010011110000101100001000110010001000100001001000110010100100101101001100000011110101001100010010010011111000111010,
	960'b010010010101010101011001010101000010110100011110000111110001110100011100000110110011000001011101010001010010111001000110010010010101011101100001010011110011101101000011010111010110101001101100011001100110001101100111011010110110110101101110011011100110101101100010010110110100111101001010010011000101001001011101011001010110111001110101011101000111010001110011011100110111001101110100011101000111010101110110011101110111011101110111011101110111100101111100011110110111101101111001011101110111011101110111011101110111011101110111011101100111010001110011011100100111001101110010011100010111001001101110011000100101100101100001011011100111001001101100010110010011110000110100001111110011111101000111010111100110000101011001011010010110111001100100011000010110101001110100011110000111100001111000011101110111100001111000011101000111001101101110011001000101010101000001001011000010001100100000001000010010001100100111001011000011010100110010001011000010110000110011,
	960'b011010100111010101100111010000100010001100100000001000010010001000100000001000000011101101101000010110100010110100110001010010110100111101011010011001000100110100111101010101000110101101101101011011000110101101101000011011000110110101101110011011100110100101100001010110010100111001001000010010010100111101011100011011010111000101110011011100110111010001110011011100110111001101110011011101010111011001111000011101110111011001110111011110010111110101111101011110100111100101111011011110010111100001111001011110010111100101110111011101010111010001110011011100100111001001110001011100100111001001110010011011000101111101010010010101010110011001101100010110110011110100101110001100010011010100111110010011000100111101010100010111000100111101001111010111010110110101110111011110000111100001111000011110000111011101110111011101100111010001110010011011010110000001001011001110000010101000100010001000010010001000101111001101010010100000100111001011010011010000111101,
	960'b100000100111110001001111001001110010000100100110001011000010010100100011001011100101110001110001011001100100001000101000001101000101001001010111011001000110011101001101010011100110101001101101011011000110101101101011011011000110110101101111011011100110110001100110010110000101001001001000010001000100110101010100011001100111000101110011011101000111010001110100011101000111010001110100011101100111011001110110011101110111101001111100011111000111111001111010011101010111100001111100011110110111101101111011011110110111101101111000011101000111001001110001011100010111001001110010011100100111001001110011011100110110111101100100010110010101010001011101010111000011110000101010001011000011001100110110010000000100110101001011001110100011111001010111011011000111011001110111011110000111100001111000011101110111011101110110011101100111010101110001011001110101111101010001010000110011000100101000001000110010011001000011001101100010010100101111010000010100101001001100,
	960'b100001010110010000101110001000000010011000110001001111100010100100100011010001100111011001111011011101110110010101000001001001010011101001011011011000010111000001100110010100110110001101101101011011000110110101101101011011010110110101101111011100000110111101101000010110000100111001000101001111110100100001010101010111110110101001101011011011010110111001101110011011100110111001101110011011110110111101110010011110001000001010000100100001011000011010000101100001101000100010001001100010011000100110001001100010001000011010000010011111010111100001110110011011110110101101101011011010110110110001101100011011000110110001100111011001010101111001001111010010100011110100101100001011000010111000110010001111000100010000110101001101010100100001011111011011110111011001110111011101110111011101110111011101110111011101110110011101100111010001101110011000010101010001001011010001000011101000101110001001110010011100110011001010010010101000110100001110110100001101001000,
	960'b011000110011100100100010001001110011001100111110010010110010111100100111011000011000001010000011100000110111111101011111001011010010100001000100011000010110110101110000011001000110000101101101011011010110111001101110011011110111000001101110011010110110100101011110001110100011010000110101001100100011001000110100001101010011001100110010001101000011010100110101001101010011010100110101001101100011001100110010010011101001001010110011101111011100100111010010110111011110001011100101111001101110010111100011110111011101000011000111101111011011000110010110010101000011001000110001001011110011000000110000001100010011001000110001001100110011001100110001001100010010111000101011001010110010110000101111001101110100101000110011001111110101001001100101011100010111010101110100011101010111010101110101011101000111010101110101011101000111001101101011010110010100010100111001001100110010101000100000000111000001111000100000001000110010110100110100001111010100110001010101,
	960'b001111010010011100100110001101100100100101010011010100100010111100110000011100111000011010000101100001101000001101110100010001100010011100101111010101000110101101110001011100010110100001101100011011100110111101110001011100010110101101011001001111010011101001000000001111000011101000111101001111010011111000111101001101110011010100110010001100110011001100110011001100110011000100110001001100110011010000110001001100010100011110001000100101011001101010011110101000101010010110100110101001111010011010100101101000111001110110011010100101011000100001001011001100000011000100110101001100100011001100110010001100110011001100110000001100000011001000110100001101000011010000110100001101010011011000111000001101100011010100110011010010100101000101010101010111100110101001110001011100100111001101110010011100010111001001110100011100100110000101000101001101010011000000101111001010110010010000011101000111000001110100011101001000000010001100101001001111010101011101100001,
	960'b001010010010011100110101010010110101111001101011010111000010111101001001100000001000010110000101100001011000010001111100011000010011001100101110010000010110100101110100011101010110110101101110011100000111000101101110011010100011110000111100001111110100010101001011010011000100110101001110010011000100100101000111010001100100100101001001010010000100011101000110010001110100010001000100010001010100010101000100010000110100001101000111010010000100100001000111010001110100011101000111010001100100011101001000010010000100100101001001010010000100011001000100010000110100010001000111010001010100011001000100010001000100010001000001010000100100001101000100010001010100010101000101010001010100001101000110010001100100010100111111001110110011011000111100001111010100110101100101011100010111000101110001011100010111001001110010011000100100000000110011001110000100011101001101001101100010101100100011001000110010001100100100001011010010100000100100001010000100000101011011,
	960'b001011000011010001001000010110100110111001111011011011110011011001100010100001011000010110000100100001011000001110000010011101110100100100110011001110010101110001110111011110000111001001110010011101010110110101000010010000010100100101011010011100001000011110011010100110111001011010001101100010111000101010001010100010001000011010000110100001011000010110000101100001101000011010000111100010011000100110001001100010001000100110001000100001111000011010000101100001001000010010000100100001001000010010000101100001011000011010000101100001011000001110000011100000111000010010000011100000101000001010000010011111101000000010000000011111110111110101111110100000011000001010000010100001001000100010010011100101101001000101110101010111010100101001000000001110100011010101001101011010110111001001110001011100100111001101100100010001100011011100111110010101100110101001011010001101110010110000100101001000110010001100101110010001010011101000110000001001110010011100110010,
	960'b001101110100101001011000011011010111100110000011011101100100000001110011100001101000010110000101100001011000010110000100100000100110000100111101001111100101010001110110011111010111100001110101011100110100110101001010010100100110110110000101100101101001010101101010010011110011111100110110001101010011010100110101001101010011001100110011001100110011010000110100001101000011001100110011001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110011001100110011001100110011001101000011001100110011001100110011001000110011001100100011001000110010001100100011001000110010001100010011001100110011001100110011010000110100001100110011011101001100011000110111111110010111100011010111011101100001010100000100100101001001011001100111000101110011011100100110011101000110001110000100001001010111011011110111000001011010001111000010101100100010001000100010001100110110010111110101111101001111010000010010111000100111,
	960'b010000100101110101101010011111001000010010000101011011010100010101111110100001111000010110000101100001011000010010000011100000100111010001010000010010000101101101110001011111110111101001011110011001010110000101111011100011100101100000101111001100000100001101011010011000000110001101100010011000010110000101100000010111100101110101011100010110100101101001011001010110010101100101011001010110100101101001011011010110110101110001011110011000000110000101100001011000100110000101100001011000110110000101100001011000010101111001011101010111000101101101011010010110100101101001011001010110010101100101011001010110110101110001011110010111100101111101100001011000100110001001100010011001000110001101100000010110110101000100110100001011100101000010000101100010010111001001110001011011010111000001110100011011000100110000111011010010100110000001110001011101110111000101100100010001110011001100100100001001000010100000111001011001110111011101110001011001100100100000110011,
	960'b010100100111001101111111100001011000100010000101010110010100110110000010100001001000000110000100100001001000010010000100100001001000000001100111010011110110100001111011011110110110011001101110011010101000000010010011011100110011000100111101010100110110000001100111011001100110011001100100011000110110001101100010011000010101111101011111010111100101110101011101010111010101110001011100010111010101110101100000010111110101111101100001011000110110010001100011011001000110010001100011011000110110001101100100011001000110000101100000010111110110000001011111010111100101110101011101010111010101110101011110010111110101111101100000011000000110001001100011011001000110010001100100011001010110010101100101011001010110001001010101010000100010110000111000100101001001010010000000100000000110110001110100010111000100000101001011011001110111011001111100011110110111100001101010010001110010110100100110001001110010111000111111011001010111111010000000011101100110011001001111,
	960'b011001111000000010000111100010001000011110000000010001010101110110000010100000101000000110000100100001101000011010000101100001011000010101111000010110010110101001111001010111100110101001111001011111001000110001100000001100110101001101100010011001010110001101100001011000000110000101100011011000110110001001100001011000100110000101100000011000000101111101011111010111110101111001011110010111100101111001011111010111110101111101100001011000100110001001100001011000100110001001100011011000010110001001100010011000100110000101100000010111110101111101011111010111100101111101011111011000000101111101011111010111110101111101100000011000010110000101100001011000100110010001100011011001000110001101011111011000000110000101100011011000110101011101000000010101111001000110001100011111110111110001100110010011110100110001101001011110110111111101111110011111000111100001100110001111000010110100110000001011000011011101001110011100011000001110000011011111010111010001100101,
	960'b011101011000010010001000100010001000100001110100001110110110111110000101100001101000011010000111100001111000011110000111100001111000011110000100011100000111000001000111011010010110011101101110010011000011111001011010011001010110001001100000011000110110010101011110010110100101101001011011010110110101101101011011010110100101101101011011010110010101100101011000010110010101101001011010010110100101101001011010010110100101101001011011010110110101110001011011010110110101101101011011010111000101101101011010010110100101101101011011010110100101101001011000010110000101101001011000010110010101100101011001010110100101101001011011010110100101101101011011010110110101110001011100010110110101101101011011010110110110000001100011011000010110000101100001010111000100000001000110100010000111101101111111011001010101101101111100100000011000000001111111011111010111101001100010001101100011010101000010001100100100001001011101011110111000010110000101100000000111100001110010,
	960'b011111101000011010001000100010011000011101100001010000000111111010001001100001111000011110001000100010001000100010001000100010001000100010001000100000010111010101001001011000000110011001110100001111000101101101101011011010000110000001100100011000010101110101011010010110100101100101011001010110010101101101011011010110110101101101011010010110100101100101011001010110010101101001011010010110010101100101011001010110010101100101011010010110100101101001011011010110100101101101011010010110110101101001011010010110110101101001011010010110010101101001011001010110100101101001011001010110100101100101011001010110010101100101011010010110100101101101011010010110010101101001011010010110010101100101011010010110110101101101011101011001000110001001100010011010000101110100111101010100001000001001110111011011100100011101110111100000101000000110000000011111110111101101011000001101100100010001010100001101110100111001101011100000101000010110000101100001000111111101111010,
	960'b100001101000011110001000100010011000010001001011010100011000011010001001100010001000100010001000100010001000100010001000100010001000100010001000011110110100001001001001011001100110110101000000011001000110100101100101011001010101111101011101010111000101101001011011010110100101101101011011010110110101101001011010010110100101100101011001010110010101101001011010010110010101101101011010010110100101101001011010010110010101100101011010010110100101101001011010010110010101101101011011010110100101100101011010010110100101100101011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011001010110100101101001011010010110100101101001011001010110100101101001011010010110010101100101011100010111100101111001100001011000110110010101101000011001000111100110001111011011110100001000111101011101111000001010000010100001000111111001001101001111110101111101110000001111100101011001110110100001001000010110000101100001011000001001111101,
	960'b100010001000100010001000100010010111101000111011011001101000100110001010100010011000100110001001100010011000100010001000100010001000100110000011001101100011010001001001011010110101000001001110011001110110011101100101011001100101111001011011010110110101101001011010010110100101101001011010010110100101101001011010010110010101100101011001010110100101101001011001010110100101101001011001010110100101100101011010010110100101101001011001010110100101101001011001010110100101100101011010010110100101101001011010010110010101101101011010010110100101101001011010010110100101100101011010010110100101100101011010010110100101101001011010010110100101101001011001010110100101100101011010010110100101101001011001010110000101100001011010010111000101111001011101011001100110010101101001011010100100110010000110100000000100001100110000010000110111111110000110100001100111100101000111010011010111010101111111010010100101110010000000100001011000010110000101100001011000010001111111,
	960'b100001111000011110001001100010010110011000111010011110101000101010001001100010011000100110001001100010011000100110001000100010011000100101111010001100110011100101001011010010000101110001101010011001010110011101100010010111100101110001011100010111000101101001011011010110010101101001011010010110010101101001011001010110100101101001011011010110010101101001011010010110100101101001011010010110010101101001011010010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011001010110010101101001011001010110100101101001011010010110010101101101011001010110100101101001011010010110100101100101011001010110100101101001011010010110100101100001011001010110100101101001011010010110100101101101011011010111000101110101011101011000000110100001100100011001100110000101001101011111010100101000101101001100000111100010000111100001100110101101000100010111000111111110000100010101010110001110000110100001101000011010000110100001101000010101111111,
	960'b100010001000100010001010100001110101001001000111100001001000101010001010100010101000101010001010100010101000101010001001100010101000001000110101001011110011111101010011010010100110101101101010011001010110010001011110010111010101110001011100010110110101101001011010010110100101101101011010010110010101101001011010010110100101101001011001010110010101100101011010010110010101101001011001010110010101101001011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101001011010010110010101100101011010010110100101101001011001010110100101101001011001010110100101101001011010010110010101101001011010010110100101101001011010010110100101101001011001010110010101101101011101010111100110000001100110011001000110101101001111011000100101010100110010001010000011100010000001100001100110001001001011011011001000011010000101010101110110000110000110100010001000011110000111100001111000010110000001,
	960'b100010001000100010001001100000010100001001011101100010001000101010001010100010101000101010001011100010101000101010001001100010101000001000110000001100010100010101011011010111100110100101100110011001100101110101011101010111000101110001011100010110110101101001011010010110100101101001011001010110100101101001011001010110100101100101011010010110100101100101011001010110100101101001011001010110100101100101011001010110000101100001011000010110010101100001011001010110010101100101011000010110000101100101011000010110010101100001011001010110010101100001011001010110010101100001011010010110010101101001011010010110100101101001011001010110100101101001011010010110100101101001011010010110100101101001011010010110110101101001011000010110010101101001011100010111010101101101100011011000100110100001100010010100000110000000111100001010000010101001111111100001000101111101011011011110001000100010000111010110100101101010000110100010001000011110001000100001111000011010000101,
	960'b100001111000100010001001011101100011101001110001100010001000100110001001100010101000101010001010100010101000100010001001100010000111101000110010001110100100110101011011011010010110001101011110010111100101110001011101010111010101100001011000010110110101101001011010010110100101101001011001010110010101101001011010010110100101101001011001010110100101101001011010010110010101100101011000010110010101100001011001010110010101100101011000010110000101100101011001010110000101100101011001010110000101100001011001010110010101100101011001010110010101100001011001010110000101100101011000010110010101100101011001010110010101101101011010010110100101101001011010010110100101100101011010010110100101101001011010010110100101101101011010010110110101110001011100010111000101101101011100011000110110001001100101010110110110100001001100001011010010111001111111100001010110101001101101100000101000101010001001011000100101001010000110100010011000100010001000100001111000011110000101,
	960'b100001101000100010001000011000100011111001111101100010011000100010001001100010011000100110001010100001111000011010001010100000010011101100101110001111110101000101010111011001010110000001011101010110100101110101011100010110110101101001011001010110110101101101011010010110100101101001011001010110100101100101011010010110010101100101011010010110100101101001011000010110010101100101011000010110010101100001011000010110010101100001011001010110010101100001011001010110010101100001011000010110000101100101011000010110010101100101011001010110010101100101011001010110000101100001011001010110010101100101011001010110010101101001011010010110010101101001011001010110100101100101011001010110010101100101011010010110110101101101011011010110110101101001011001010111010101101101011011010111110101111101100100011001000110011101010000001100110010111110000001100001100111101010000000100010001000101010001010011010100100110010000101100010101000100110001001100010011000100010000110,
	960'b100001101000100010000110010011010100101110000100100010001000100010001000100010011000100110001001100001101000100010001001011111100010011000110010010001010101011001011100011000000101111001100010010110110101110001011011010110110101101101011010010110110101101001011010010110100101101001011010010110010101101001011010010110010101101001011010010110100101101001011010010110010101100101011001010110010101100001011000010110010101100001011000010110000101100101011010010110000101100101011001010110010101101001011001010110010101100101011001010110000101100101011000010110000101100101011000010110010101100101011001010110000101101001011001010110100101101001011010010110010101101001011010010110010101101001011010010110100101101001011001010110100101100101011010010110100101101101011011010110110101110001100010011010000110001101010011001111000011010010000001100010011000010010001001100010111000101110001011011100000100010010000010100011001000101010001001100010011000101010001001,
	960'b100001011000100101111101001110100101111010000101100001111000011010000110100001101000011110001000100001011000100110001011100000000010010100110101010001010101100101100001011000010101111001100100010111010101101101011011010110110101101001011011010110100101100101011010010110100101100101011010010110010101101001011001010110010101100101011001010110100101101001011001010110010101100101011001010110010101100101011000010110000101100001011001010110010101100101011010010110010101100001011010010110000101100101011000010110000101100001011000010110000101101001011000010110010101100101011000010110010101100101011000010110010101100101011001010110110101101001011001010110010101101001011010010110100101101101011011010110100101101101011011010110110101100001011010010110110101101101011011010110100101110101100001011001110101111101010000001111010011011110000010100010111000101010001010100010111000101110001100011101110100000001111101100011001000101010001001100010101000101010001010,
	960'b100001101000100001101011001101000110111110000011100000111000010010000100100000101000010010000101100001011000100110001011011111110010010100110111010001110101110001100101011000100110000001100011010111010101110101011011010111000101101001011010010110100101101001011010010110010101101001011001010110010101101001011010010110010101101001011010010110100101101001011000010110000101100101011000010110100101101001011001010110010101100101011001010110110101100101011000010110010101100001011001010110000101100101011001010110000101100101011001010110000101100101011001010110000101100101011000010110100101100001010111010110100101100101011011010110100101101001011010010110010101100101011010010110100101101001011010010110100101101001011010010110100101100001011010010111000101110001011100010110110101111101100010011001110101111001001101001111110011101110000011100010111000101010001010100010101000101010001011011110110011110101110110100011001000101010001010100010101000101010001010,
	960'b100001101000010001010001001111000111110010000100100000101000001110000010100000101000001010000001100000111000001101111001011001110010011100111110010001110101111001110000011010000110001101100110010111010101110001011101010111000101101001011010010110100101101001011010010110110101100101011010010110010101101001011010010110010101101001011001010110100101101001011010010110010101100001011001010110000101100001011001010110000101100001011000010110000101100101011001010110010101100101011001010110000101100001011001010110010101100101011001010110000101100101011001010110010101100101011000010110010101100101011000010110100101101001011010010110100101100101011010010110010101101001011010010110100101100101011010010110110101101001011010010110100101101001011100010111000101101101011100010111000110000101100101011010100110000001001000010000110100000010000100100011001000101010001010100010101000101010001011011111100100000001101111100011001000101110001011100010111000101110001011,
	960'b100010000111111100111100010011111000001110000101100000111000010010000100100000111000001101111111100000000111011001110000011010010010101001000010010001110101101101110001011010100110001101100101010111110101110101011110010111000101101101011000010110110101101101011001010110110101101001011010010110010101100101011010010110100101101001011010010110010101100101011010010110010101101001011010010101110101100001011000010110010101100001011000010110000101101001011001010110000101100101011001010110010101100001011001010110100101100101011001010110000101100001011001010110010101100101011000010110010101100001011001010110010101101101011010010110100101100101011001010110100101100101011010010110010101100101011010010110100101101101011010010110100101101101011011010111000101110001011110010111010110001001100111011011000101110001000110010001100100001110000100100010111000101010001010100010101000101010001011100000110100010001100110100011001000110010001011100011001000101110001011,
	960'b100011010111010100110010011001101000011010000110100001001000001010000011100000101000000101111100011110110111011001111101011101010010110001001100010001100101001101110011011011010110011101100110011000000101111001011110010111010101110001011011010110100101101001011010010110010101101001011010010110010101101001011001010110010101100101011010010110010101100101011010010110010101100101011001010110100101101001011001010110100101101001011001010110100101100101011001010110010101101001011001010110010101100101011001010110010101100101011010010110010101101001011001010110010101101001011010010110100101101001011010010110100101101001011010010110010101101001011001010110010101100101011001010110100101101001011011010110100101101001011010010110010101110001011100010111100101110001011111011000010110010001101011011100010101001101000100010100000100100110000101100010111000101010001010100010101000101010001011100001100100101101011011100010111000110110001100100011001000110010001100,
	960'b100011100110000000110011011101111000011110000110100001001000000010000010100000010111111101111010011111010111110101111110011101110011000101010101010011010100110101110000011011110110100101100101011000010101111101011110010111000101110001011100010110110101101001011010010110100101100101011010010110010101101001011001010110100101101001011001010110100101101001011010010110010101101001011010010110010101101001011010010110100101101001011010010110100101101001011011010110100101101001011011010110110101101001011011010110100101100101011010010110110101101001011010010110100101101001011001010110010101101001011010010110010101100101011010010110100101100101011010010110100101101001011010010110100101101001011011010110100101101001011011010110010101110101011100010111110101110101011111011001010110011101101110011100100100110101000110010110100100111010000100100011001000101010001010100010101000101010001011100010000101001101001111100010011000110010001011100010111000110010001011,
	960'b100010000100010001000001100000111000011110000111100001000111111010000010100000100111110101111010011111100111111001111111011101110011011001100001010111010100100101100101011100010110101001100110011000110110000001011110010111100101110001011100010110010101101001011010010110100101101001011010010110010101101001011010010110010101101001011010010110100101101001011010010110100101101101011010010110100101101001011010010110100101101001011011010110100101101101011011010110110101101001011011010111000101110001011011010110100101101101011010010110100101101101011011010110100101101001011001010110100101101001011010010110100101100101011001010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101110001011100010111100101111101100010011010010110101101110001011101100100100101001110011000110101010010000101100010111000101010001010100010011000101010001011100010010101111001000011100001001000110010001011100010111000101110001011,
	960'b011101010010111101011001100010101000101010001001100001110111111010000010100000100111110001111011011111110111111110000000011100100011111001101100100000100100110001001101011101110111000101101010011010010110001001011111010111010101110101011100010110100101101101011010010110100101101001011010010110100101101001011001010110100101100101011001010110100101101101011010010110100101101101011010010110100101101101011011010110110101110001011100010111000101110001011101010111000101110101011101010110110101101101011011010111010101110001011100010111000101101101011011010110110101101001011011010110100101101001011011010110010101101001011010010110100101101001011001010110100101101001011010010110100101101001011010010110100101101001011010010111000101110001011011010111110110000001100110011010110110110101111001011101000100011001110011011100100110000010000100100010011000100110001001100010001000100010001010100010100110101000111010011111001000110010001010100010101000101010001010,
	960'b010101010010101101101100100001011000010010000100100000100111100101111110011111100111010101111000011110100111101001111011011011000100010101101010100010010110001001000111011101110111010101101100011010100110010001100000010111010101101101011011010110110101101101011010010110100101101001011010010110100101101101011010010110100101100101011010010110100101101001011011010110100101101001011011010111000101110001011100010111000101110101011101010111100101111001011101010111010101111001011110010111100101111001011101010111010101101101011101010111010101110001011011010110110101101001011010010110100101101001011010010110100101101001011010010110010101101001011010010110100101100101011010010110100101101001011010010110100101101101011011010111000101110001011100010111100110001001101000011010000111000101111011011001110101010110000101011101000110010010000100100010001000100010000111100010001000100010001000100010100111010000111000011100111000101110001010100010011000100110001001,
	960'b001100010011101001000111010010100100101001001010010010100100100101001001010010010100100001001001010010010100100101001001010010010101111101100010011111011000101101011001011000010111011101110000011001100110011101100110010111010101101001011011010111000101101101011001010110100101101101011011010111000101101101011010010110110101101101011011010110110101101101011011010111000101110101011101010110110101110001011101010111000101110101011110010111100101111001011110010111110101111001011110010111100101110101011101010111010101110001011101010111010101110001011101010111010101110001011100010110110101101001011010010110100101101101011011010110100101101101011011010110110101101101011010010110110101101101011011010110100101101001011011010111000101101001011100011000010110100001100101011010100111011101101011010011101000010110000110011011010101111010000011100010001000011110000111100010001000100010001001100010100111101100111011011001011000100110001001100010001000100010001001,
	960'b001000010101100001000111010010110100101101001011010010110100110001001100010010110100101101001011010010110100101101001011010001110110111101011110011010010111111101110011010011100110111001110101011001100110001001100111011000010101110101011100010111000101110001011100010111010101110001011011010110100101101101011010010110110101101101011011010110010101101101011100010111000101110101011110010111000101110101011101010111010101110101011101010111100101111101011101010111110110000001011110010111010101110101011101010111000101110001011101010111010101110101011100010111000101110101011101010111010101110001011100010110010101101001011011010110110101101101011010010110110101101101011011010110110101101101011100010111000101110001011100010111010101101001011011011001100110010001100110011011010111001101010011010000111000110001111011011001010100111010000001100001111000011010000110100001111000100010001000100010101000000001000010010110001000011110001001100001111000011110001000,
	960'b001001110101000101000111010011000100010101000011010000110100001101000011010001000100011101001000010010010100010101001011010010010111000101001010010100110110011001110011010001100101011101110010011010100110001101100010011001000101111001011101010110100101110001011101010111000101110001011011010110110101101101011010010110100101101001011010010110100101101101011100010111000101110101011110010111000101111001011110010111100101111101100000010111110101111101100000010111110110000101100000010111110110000001100000010111110101111001011110010111010101110101011111010111010101111001011101010110110101110001011100010110100101101101011011010110100101101001011010010110110101101101011011010111000101101101011100010110110101110001011100010111000101101101011011011000010110001001101000011011110110000001000100010001110111101001100111010111000111101110000100100001001000010010000100100001011000010110000101100001101000001101001110010011011000010010001001100001111000011110001000,
	960'b001010010011010001000011010011010100001100111000001110000011100100111000001111010101110101100111011011000100100001001011010010100110101000100101001110000100010001001001010010100011111101001100011011110110101101100100011000010110010001100010010111100101110101011111010111100101110101011101010111010101110001011100010111010101110101011101010111010101111001011110010111010101111001011111011000000101111101100010011000010110001101100011011000110110001101100100011000110110010001100011011001000110001001100011011001000110001001100010011000100110000001011111010111100101111001011101010111010101110101011101010111000101110101011100010111010101110101011110010111010101110101011101010111100101111001011101010111000101110001011011010111110110010001100000011000110110011101101111011010110100001101001010011001110101001101000111001010110111110010000110100001011000010110000101100001011000010110000101100001101000010001011011010001101000000010001000100001111000100010001000,
	960'b001010110011000101000011010011010100001100111010001110010011011100110101001101110011111100111110010001000100010001001100010010000111000001100101001000110011011000111001010010010011111001000010011001110110111001101000011001000110000001100100011001110110001101011111010111110101111101100000011000000101111101011111011000000101111001011111010111100101111001011110010111110110000001100001011000100110001001100011011000110110010001100101011001010110010101100101011001100110011001100101011001010110010001100101011001010110010101100010011001000110001101100010011000100110000101100000010111100101110101011101010111000101110001011100010111010101110101011111010111110110000001100000010111110101111101011101010111000101110101100010011001000101111101011111011001110110101001101011010101100100000001010101010100110100000100110010011101011000011010000110100001101000011010000110100001011000010110000110100001111000011001101011010000000111100010001000100001111000100010001000,
	960'b001011100011000101000011010011010100001100110100001101100011100000110100001100010011000000110001001100100100001101001100010010000110111101110001010000110001000000101000001100010011010000111100010000100100110101100110011011100110101001101000011001110110010101100110011010000110100101101010011010010110101101101010011001110110100001100110011001110110011101101000011010000110011101101000011010100110101001101011011010100110101101101011011011000110110001101011011011000110110001101011011011010110101101101011011010110110101101101010011010010110101001101001011010010110100101101010011010000110100001100111011001110110100001101000011001110110011101101001011010010110101001101001011010010110101001101001011010000110010001100101011001010110011101101100011011010101100101000100001111010100010101000010001110000001100000101010100000001000100010000110100001111000011110000111100001101000011010000110100001101000011101110110001111100110110010001000100010001000100010001000,
	960'b001011100011000101000011010011010100001000110010001100010011000100101100001010000010011100101001001011100100001001001100010010000110110001110000011001110001111100010100001001010010111100110000001101000011111001001010011000000110111001101101011011000110110001101010011010010110100101101001011010000110101001101001011001110110011101100111011001110110011001100110011010000110100001101000011001110110100001101010011010010110100101101010011010100110101001101011011010100110101001101011011010110110101101101010011010100110100101101010011010000110100001101001011001110110100001101000011001110110100001100111011001100110011101100111011001110110011101101001011010000110100101101010011010010110101001101001011010010110101001101101011011010110101001101101010101100100000000111001010000010011111100111001001011000001100101110110100010011000100010001000100010001000011110001000100001111000011110000111100001111000100101111111010000000101110010000111100010011000100010001001,
	960'b001011110011000001000010010011010100001000110010001100100011000000101001001001010010010100100111001010110100001001001100010001100101010001010011011001010110001100111011000110010010011000100110001011000011001100111001001111010100101101011101011011100111100001111101011111010111101101111000011101110111011101110101011100110111001101110001011100100111000101110001011100010111001001110011011101000111001101110101011101110111011101110110011101110111100001110101011101110111011101110101011101110111011101110101011101000111010101110101011101000111010101110011011100100111001001110100011100100111000101110000011100000111000001110001011100010111001101110110011101100111100001111001011110000111100001111000011110010111101110000000011011110101001101000100010001100100011000111100001110100011010100100110000111100111011110001100100010101000101010001010100010011000100110001001100010011000100110001001100010011000101010000100010010010100111110000110100010101000101010001010,
	960'b001011110011000001000010010011010100001100110001001100000011001000110001001011000010101100101011001011100100001001001101010000110011011000110010010000000101010001001110000100000001011000101010001010000010101100110010001111000011111001000001010010100101101001110101100000001000001010000101100001001000010110000011100000101000001010000000100000011000001010000011100000101000010010000100100001101000011110000111100001111000100010000101100010001000100010000110100001011000011010000110100001011000010110000111100001111000011010000110100001101000011110000101100001011000010010000010100000011000001010000010100000001000000110000010100000101000010010000101100001101000100010001000100001111000011010000100100000100111011101010100010001000100000001000111010001010011110000110111001100110010010100010011011110001000111010001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000110010001001010110010100001110000001100011001000101110001011,
	960'b001010110010111001000010010011010100001000110000001011100011000100110011001101010011001100110011001100110100001101001101010000110011001100110000001100000011100000111111001110010001000000010110001001010010011100101100001100100100001101000010001111010011111001001001010101010101111101101100011100000111000001110010011101110111011101111000011111011000000110000010100001011000100010001001100010111000110010001111100100001001000110010010100100111001001110010011100100111001001110010100100100111001001010010001100100011000111110010000100011111000111010001011100010111000101110000111100001101000011010000101100000011000000001111111011111010111101001111001011110000111010101110100011100010110110001011100010100010100010101000000010010000101001101001100001110100011001100101101001100010001010100011001100001101001000010001110100011111000111110001110100011101000111010001110100011011000110110001101100011011000110110001101011010100011110001111001100011101000110010001100,
	960'b001010000010110001000010010011010100001000110001001100000011000100110010001100100011000100110100001100110100001001001101010000110011001000110010001100100011011100111001010001000100001100011101000011000001110000101110001011110011000000110000001100010011010000111111010010000100111101001110010011100100111001001111010011100100111001001101010010100100101001001011010010110100100101001010010011000100111001010000010101010101100101011101010111100110000001100001011000110110001101100101011001000110010001100011011000110110000001011101010110110101011101010110010101010101001001001111010011010100101001000111010001000100010101000101010001010100010101001001010011000100110101001110010011010100111001001101010011010100001100110110001101000011011100110010001101000010011100001101000111010111110110001000100100001001000110010001100100011001000110010000100100011001000010010001100100011001000010010000100100001000111110010000011110000011100101101011100011111000111110001101,
	960'b001010010010101001000010010011010100010101000011010000100100001001000010010000100100001001000011010000110100010101001100010000100011001000110011001101110011011100110111010000110100101001000111000011110000110000010001001000110011000000101011001010110010111100110100001101100011100000111010001110110011101000111001001101000011001000110000001100010011000000110000001011110010111000110000001100100011010000110100001101100011100100111100001111000011111001000000010000100100001001000010010000000100000001000000001111100011110100111100001110110011100100110110001101100011010000110011001100010011000000101111001011110011000100110010001100000011000100110011001101010011100000111000001101110011100000110111001110110011100000101111001010100010111000110001000101110001001100011010011111101001010110010101100101001001010010010011100100111001001110010011100100111001001110010011100100111001001110010011100100101001001010010011100000110011110001011001100011111001000110001111,
	960'b001010100010110001000010010011000100110001001101010011010100110101001101010011010100110101001101010011010100110101001100010000110011001100110001001101100011010100110100001111100100100001001100010010110100001100100001000011110000100100010001001001010011111001010001010011100100100001000110010001110100011101000111010001000100001101000101010001100100010001000011010000100100000101000011010000110100010001000110010001110100011101001001010011000100110101010000010100010101001001010001010011110101000001010000010011110100110001001001010010010100100001000111010010000100011001000110010001010100011001000101010001010100011101001000010010100100110001001010010010100100111001001101010011010100110001001111010101110101101100111111000111010000110100001010001000011000000110001101100101101001011010010110100101101001011010010110100101101001010110010101100101011001010110010110100101101001011010010110100101011001010110010101100011000100010101001010100011011001001010010001,
	960'b001010100010111001000000010000110100001101000011010000110100001101000011010000110100001101000011010000100100001001000010010000000011010000110011001100100011000100110111001111000100001101000111010010000100110001001100010010100001010000001001000010010001000100101011001110110100010001010111010011010100010001000110010101000101000101000100010000010100000000111111010000000100010000111101001111010011111001000001010000110100011101010010010010100100110001001110010100110101010001010101010111100101001101001111010011000100100101000111010001100100111101000110010000110100001000111111001111100100000101001100010000010100000001000001010000110100010101010100010100010100010101000101010011100101010101000011001111100010110100001101000011110000100000011111100001101001101110011011100110001001100010011001100110001001100110011001100110001001011110010111100110001001100010011000100110001001100010010111100110001001011110010111100100110101010000111111100001111001010010010010,
	960'b001010010010110100110010001101100011100000111001001110010011100000110111001101100011001000111000001011110010111100110001001100010011001100110101001011110011001100111001001110100100000001000001001111000100000001000011010001110100111100101011000100100000110000001100000011000001101110011011010101000000111100011010100010111000000100011110000100010001001100010101001101010101110000011010000101000001010100010110000101010011000101101111000111100001010100011000000110100001100000101100011111010010011100011000000110000001100100011000001001110111101100101100000110000001100100011000000101110010010101111010001010110001011000011000000110000010110010010010100001100001111100010011011001011001111100100011000101010001001000011101011111110101011010001011100111101001110010011100100111001001101110011100100111001001101110011001100110001001101010011001100110011001101010011010100110101001101010011001100110011001100110011001100110000110100000111100100000001001011110010101,
	960'b001010100010110000101111001100100011011000111001001110000011100000111000001101000011010100111001001011100010111100110011001100110011010000110101001011100011001000110110001101100011101000111111001111100011111000111001001101010011110101000011010001000100001000111011001110100100000101001101001111110011100101000011010100010101010101010000010101010101111101100010011001010110110001100111011001010110010101100100011000100110011001101111011001100110100001101011011011000110110001110010011111000111011001110111011110010111101001111010011111111000100001111110011111000111101101111100011110110111111110001001100000010111111110000000100000011000010010010010100101011000011001000100011000011001110110010010100100011001000010010011101000011001111010100100101000111010001010100010101000111010010010100101101001011010011010100101101001011010010110100101101001001010010110100100101001001010010010100011101000111010001010100010101000010111100100110111011110101010000010011110,
	960'b001100010011001100110101001101100011011100111010001110110011110100111110001111010011111101000010001111010011110101000001010000110100001001000010001110100011011100110111001111010100001101000111010001000100011101001010010010100100101001001100010010110100110001001100010011100101000001010000010101010101011001010101010101010101110101100101011011010111001101110011011100100111000101110011011100110111011001110111011101110111100001111000011110110111111110000001100000111000001110000110100010001000110110001111100111011010000010010101100101101001010110010110100101111001011010010110100101101001100010011000100110111001110110011110101000011010001010100010101010001010011101011000010110101010011010101100101010101010101110101011101010111010101110101010101010101010101010101010101010111010110010101100101011011010110110101101101011011010110110101100101010111010110010101011101010111010101010101010101010011010100010100111101001011000011100111000011011101010010110100100,
	960'b001111000100000001000011010000100100001101000101010001110100011001000110010001100100011001000111010001110100100001001011010011000100110101001100010010010100100101001001010010110100101001001101010011100100111001010011010101100101010101010101010101110101101001011010010111100110010101100111011010100110101101101011011010110110110101101110011100010111001101110010011100010111000101110001011100110111011101111001011111010111111110000010100001011000010110001000100010101000101110010001100101111001110010011100101111011100001110100101101000101010010110100101101001001010001110011111101000101010001110100011101001001010010110100110101001101010100010101011101011101010110101100011010100001010100110101110101011001010110110101100101011001010101110101011101010111010110010101101101011011010110110101101101011001010110010101100101010111010101110101011101010101010101110101101101011011010110110101110101011011010110110101100101010101001011001000000011000001010100010101011,
	960'b010001010100100001001011010100000101000001010001010100010101000001010000010100000101000001001110010011000100110101001111010100000101000001010010010100100101010001010111010110100101100101010111010101100101100101011011010111100110001001100100011010100110110101101100011011000111000001110010011100100111001001110011011101000111010101110110011101110111100001111000011110000111100001111001011111011000001010000111100100001001010010011100100111001001000110010001100100011001000110011000100111001001110010011111110000011100101110101010101001111010100010100111101001111010011110100110101001111010010110100101101001011010011010100110101000111010011110101010101010111010101101101111010000101010010010101011101010011010100010100111101010001010101010101010101010111010111010110010101100001010111110101110101011001010110010101101101011011010110010101011101010101010101010101010101010111010110010101101101011101010111110101110101100001010010001001100010101101010110010110100,
	960'b010101010101010101010111010110110101110101011101010111100110000001100000011000010110000101100000010111110110000001100001011000100110001001100010011000110110001001100010011001000110010001100100011001000110011001100111011010100110110101101111011100100111001101110011011100110111001101110011011101000111010101110110011101110111100101111011011111100111111101111111011111100111110101111100011111100111101110000111100110101010010010110011101101011010111010101100101001111010001010011111100111111001111010100010101111101100001110101001101001111010011110100010101000101010001110100110101001101010010010100100101001011010010110100110101001111010100010101010101010111010110001111110001110111001100110101100101010001010100010100111101001101010011010100101101000111001101010011100101001001010001010011010100110011010000010100001101000001010010110100100101000111010010010101010101011001010110110101110101011001010100110101101101011011010011101011000010010001010010010110010,
	960'b011001100110010101100101011010000110100101100110011001100110101101101100011011010110110101101101011011010110111001101111011011100110111101101111011011100110110101101101011011100110111001101111011100000111000001110001011100110111001101110101011101100111011001110101011101100111011001110111011110000111100101111001011111101000010010001001100010111000100110000001011111010111110001111001011110100111110010001001100111011010110010110110101110001011011110110110101101011011001110110001101100001011001010110111101111011011101010110001101011111011001010110101101101001011000110101110101010101010011010100110101001101010011010100111101001111010011110100111101010001010100110000110001110001001000110101011101010011010100010101001101001111010011110100101101000101001000010000111100001111000010010000001100000001000001010000010100000011000010010000010100000011000000110001100100100101001000110001110100010011000100010001110100100101001010001011011001110111000111110100100,
	960'b011100100111001101110011011100110111001101110010011100100111001101110011011100110111001001110010011100010111000101110001011100000111000001110000011100010111001001110010011100100111001101110100011101010111010101110110011101100111011101111001011110100111110001111110011111111000000110000010100000111000010010000101100001101000011110000010011111100111101001111010011110100111101101111011011110110111101101111110100001111001010110100000101010011010101110100111101001111010101110101010101010001010101110101101101010111010101010101011101010111010111110110010101100011011001010110000101011101010110010101100101010111010110110101110101011001010101110101100101011001010110110010011001110111000101110101111101011011010101110101101101010111010110110110010101011011010001010011100100111011001101010011010100101001000111110001011100001111000010010000000011111110111111001111110100000000111111101111110011111100111110101111010011110100111100101010101001100010111000010000111,
	960'b011011100110111101110001011100110111010001110101011101100111011001110110011101110111011001110100011101000111001101110011011100110111001101110011011101000111010101110101011101100111011101111000011110110111101101111100011111011000001110001000100010101000110110001011100001011000001010000010100000011000001001111100011111000111110101111011011110000111010001110110011101110111100001111010011110110111101101111010011111011000000010000000100001001000100110001000100010101001001010011110100111001001011010011000101000011010000010011100100111101010001010100100101000111010010110100100101001011010010110100110101010011010110010101110101011111011000110110011101100111011010010100000010000110111111010100110101001011010010010100100101001101010101110110000101011111010101010100111101010011010011010101000101010011010100110100010100101111001011010010101100101101001100110010111100110011001011110010110100101111001100010010111100100011000100001100011001011110111000010010000,
	960'b011011010110110101101110011011110110111101110000011100010111001101110001011011000110101001101010011010010110100101101100011011010110110101101110011011100111000001110011011110000111110001111100011110100111010101110110100010001001110110100001100111111001111010011010100011111000001001111101011111011000000001111010011110000111010001110100011100110111000101110010011100110111010101110110011101110111100101111000011101110111100001111010011110010111101101111110100000001000001010001011100011011000101110001110101000111010000010010011100101001001100110011111100111101001110110011100100111011001110110011101100111101010000010100010101001001010011010101010101010111010101110011100010001110110101010011001100110001001011110010111100101111001101110100000100111111001110010011000100101111001100110011001100110101001101010010111100100111001001010010001100100111001010110010111100110011001100110011010100110111001110110011101100110011001011001110100001011110110011110010011,
	960'b011011100110111101101111011100000111000001110000011100000111000001101101011001000101110001011000010101100101010001010110010110000101101001011111011000010110001001101001011101111000000110000010011111010111010101111001100101101010010110101000101001111010010110100001100100010111010001101101011011100111010001110010011101100111010101110101011101000111000101110001011100100111001101110100011101100111011101110110011101110111110110000001100000001000001110000110100001011000010010001000100011001000111010010101101110011011010110011001100110011001110010100000101000001001110110011100100110111001101110011000100101101001001010010001100100101001001110010110100110001001100010010000010010100101110110010001100100011000111010001101100011001000110110001110100011101000110010001001100010011000110010010000100100101001000110001110100011001000110010001100100011001000111010010011100101001001010010010100100101001001010010010100100100111001001101111000001100000101110010010000,
	960'b011011000110111001101111011011110110111101110000011100010111000101110000011100010111000001101100011001100101101001010100010101000101011001011011010111100110001101101101011111001000101010010010100100111001001010010100100110101001100010010111100110011001110010011101100101010111111001110110011110011000000110000001100001001000001110000010011111000111011101110101011101100111011001110101011101010111011001110111011110000111110101111111100000000111111110000000100000101000010110001010100100011001010110011100110000011011111010011010100101101001010110010110100110001001100110011011100111111001111110011010100101101001000110010000100011011000101110001100100011001000101010000110010011000101001010001000100010001000001110000001100000000111111101111110011111010111110001111011011111000111110110000001100000111000011010000101100001011000010010000101100001111000101010001100100011011000111010001111100011111000111110001110100011011000111001110110001011110101001110001011,
	960'b011010110110110001101100011011000110110001101100011011000110110001101100011011010110111001101101011010010110010001100000010111100101101001011010010111000110010001110010011110111000001010001000100010111000100010000110100010011001000010011000100111001001111010100001101000101001110110011010100110101001111110100000100111111010000010100001100110111001011110010001100011111000111010001011100001111000010010000011100000011000001010000010100000010111111110000000100001001000100110001110100101001001011110011110110000011011111110011111100110101001100110011001100110011001101010011110100111111001111110011111100111101001110110011010100101101001001110010010100100011001000010001001010100110100011110000100100001010111110101111100011111000111100001110101011100110111000001101111011011110111000101110001011100110111011001111000011110000111011001111000011110100111111001111110100000011000010110000110100001111000011110000111100001101000011101110001001011000100110010000011,
	960'b011011000110110101101100011011000110110001101011011011000110101101101001011010010110100101101010011011000110110001101110011011100110110001101011011010110110100101100111011001000110001101100011011010000110100101101000011011010111100001111111100001101000101110010001100101011001100110011100101000001010001110100101101010001010101110101011101010101010100010101001101010101010100110100101100111101001110010011101100110101001101110011100100110011000111110001001100010101000111110010100100110001001110110100100110010001100010110100010100111001001101110011011100110101001100110011011100110111001110010011110101000111010010010100001101000001010001110100010100111111001110110011000011000010100001010001001100011111000101110000110100000100111111001111001011101000110111101101101011011100110111101101111011011100110111101110000011100000110101101101010011010100110110101110000011101000111011101111001011110100111101101111100011111010111110101101010001011000100100001111101,
	960'b011010110110101101101100011011010110110101101101011011010110110101101101011011010110110001101101011011100110111001101111011011110110111001101101011011100110111101101110011011010110110001101010011010010110011001100010010111110110000001100001011000010110011001101110011101100111111010000110100011111001101010100110101100001011001010110000101011001010100010100100101000111010010010100111101001001010001110100011101001001010011010100110101010001010010010100000100111001001110110100001101001011010100010101101110011001100011110100011100111101001110110011100100111001001110010011101100111111010000010100001101000011010000010011111100111111010000010100010101000011010000110100001011100010011111010010010101000001001110010011001100101101001010110010001100010011000011010000100100000101000001010000001011111110111111001111101011110100111010101110000011011100110110101101101011010110110101001101010011010100110110001101101011100100111010001100010001010110100001101110111,
	960'b011010100110101001101011011010110110110001101100011011010110110101101101011011010110110101101110011100000111000101110001011100010111000001101110011011100110111001101111011011110110111101101111011100000110111101101111011100000110111001101100011001010101110101011101011000100110010001101011011011110111011010000010100101001010001010101100101100011011010010110010101011011010101010101011101011011010011010100011101000111010001010100010101001011010011010100111101001111010010010100100101010001010100110101100110000101011110110101001101001011010010010100011101000111010001110100011101001001010010010100100101000101010000110100001101000011010001010100010101000101010000110100001011110110011110010010001101000101001110010011010100110111001111010011100100110011001100010011011100110001001000110001111100011101000111010001000011111110111101101111101011111100111110001111001011101010111001001110001011011010110100101101001011010010110101101011100001010100011111001101111,
	960'b011001100110011101101000011010010110101001101011011011000110101101101100011011000110110001101100011011000110110101101101011011010110111001101110011011110110111001101111011011110110111101110000011100000110111101101111011100000111000101110001011100010111000001101111011011010110100101100111011001000110010101100101011001100110110101110111011111101000100110010100100110011001011010010111100110111001101110011110101000101010001110100100101000101010001010100010101000011001111110011110100111111010000010100010101010011010110010101001101010001010100010101000101010011010100110100101101001011010100010101001101001101010001110100010101001001010010010100011101000111010011010101000100010000011110010010000101010101010011010100100101001001010011010100011101000011010000110011111100111101001101010010111100101011001001010010001100011001000100110000111100010001000011010000010100000001000000110000000011111100111101101110110011101000111010101100101001010110011111001110110,
	960'b010111100110001101100100011000110110001101100100011001000110010001101000011010010110100101101001011010100110101001101011011010110110110001101100011011010110110101101110011011100110111101101111011011110110111101101111011100000111000001110001011100000111000001110000011011110110111001101101011011010110110101101100011010010110011101100110011001100110101101110110100011011001010110010100100110111001110010011010100101111001011010010111100110011001111010100000100111011001110010011011100110101001101010011101100111101010000110100011101001011010010110100110101001111010100010101010101010001010011010101001101010111010100010100111101010001010100110101000101010001010011010101001100011110011100110000110101010101010011110100101101001011010011010100110101001011010001010100000100111111010000110011110100111101001110110011100100110101001011110010100100011101000110010001010100010001000100110001010100010111000100110001001100010001000100001110001001010110100000010000010,
	960'b010111000101111001011101010101000101011001011011010111010110000101100011011000110110001001100010011001000110011001100111011010000110100001101001011010100110101101101011011011010110111001101111011100000110111101101111011011110110111101101111011011110110111101101110011011100110110001101011011010100110101001101001011010010110100001100110011001010110011101110011100001011000110110010000100110001001110010011101100111011001110110011101100111011001111010011111100111101001111010011101100111001001101110011100100111011001111110100010101001101010011010100000100111101010000110100100101001001010001110100011101000111010000110100010101000111010010110100101101001111010010110100101100100010011100101111011101010011010100110100110101001111010100110101010101010011010100010101000101010001010100010100101101000101010000010011100100110001001010110010101100101001001011010010101100100111001011010010110100101001001000110010000100100001001000001111000001011010100000110000011,
	960'b011000000110000001011111010111110110000001100000010111100110000101100011011000010101110101011101011000100110010001100101011001100110011001100101011001010110010101100110011001110110100001101010011010110110101101101011011011000110110001101011011011000110101101101011011010110110101101101010011010010110011101100101011001000110001101100010011000110110011001101101011100100111010101111001100000011000011110001101100100101001100110011100100110111001101110011011100110111001101110011100100111111010000010100000101000001010000010100000101000111010001110011101100111001001110110011110100111111001110110011011100110101001100110011011100111111010001110011111100111011001111010100000100100010011111001101011100111101001110110011010100111001010010010100111101010001010100010100111101000101001111010011111100111001001110010011111101000001001110110011101100110111001101010010111100110111010000010100000100111111010000010011111100111001001101001111100001011000100001110000101,
	960'b011000000101111101011101010111110110000001100010011000100110001101100101011001010110010101100101011001100110011101100111011010000110100001100111011001100110010101100100011000110110010001100100011001010110100001101000011010100110101001101001011010010110100101101001011010100110101001101010011010000110010001100010011000110110101001110010011110000111110110000101100010101000110010001110100100011001010010010110100101111001100110011100100111001001110010011101100111001001110110011101100111101001111110011111100111111001111110011111100111111001111110011111100111111010000010100001101000111010000010011010100101111001010110010100100101011001011110010111100101101001100010011001100011000011110101011100100101001001011010010110100110001001110110011110100111111001111010011101100111101010000010100000100111101001110110011110101000001010001010100010101000111010010110100011101000111010001010100011101000111010001110100011101000111010000101111110001001110100000110001000,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = r_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		g_data = g_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		b_data = b_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		// r_data = {8{picture[(y_cnt - y_pin)][((x_cnt - x_pin))]}};
		// g_data = {8{picture[(y_cnt - y_pin) + Y_WIDTH][((x_cnt - x_pin))]}};
		// b_data = {8{picture[(y_cnt - y_pin) + (Y_WIDTH << 1)][((x_cnt - x_pin))]}};
		// r_data = 8'b0;
		// g_data = 8'b0;
		// b_data = 8'b0;
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule