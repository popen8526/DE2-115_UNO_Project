module blue_skip(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111111111111111111100111101000001001110010110111101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110001001110110100110111100111111111111111111,
	240'b111111111111011010111011110011011110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011010000110000011111011011111111,
	240'b111111011100010111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100010011111101,
	240'b110010101101001011111111111101011011010110010101100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010011100100001000111110010001100101011011010011110100111111111101001111001010,
	240'b100111111111000011111110100111100100111101010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100010100111001010110011110001000010001100111010011010100111010011011111111101111010110011011,
	240'b101011101111111011101110011001100101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110100011001011111100111111001011101111100111000101000101100100111010111111111010101100,
	240'b101101101111111111100100011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101111100011111111111101010010111000110101111111101101000010001011011111000101111111010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011110011110111111011110110111110110101001001110110001001100100101011111111000011111111010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100101011101111101101110110101111101110001011111100100111101111001101001111000001111111010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100011001110100001100000011001111110001111001010101011111101100001100110111000001111111010111000,
	240'b101101101111111111100100011000010101001101010011010100000101000001010000010011110101000001010010010101000101010101010101010101010101010101010010011010001110110010101000010011110111000111101000111111101010110101011100111000011111111010111000,
	240'b101101101111111111100100011000010100111101100000100010111010010010100011100110011000100001110001010110110101000101010001010101000101010101010101010100101001101111110111110010111011001011110000110111100110010101011110111000101111111010111000,
	240'b101101101111111111100100010111010111011011011000111111101111111111111111111111111111110111110010110110001010111001111010010101100101000101010101010101000101010110001110110011111101110010110101011010100101000001100000111000101111111010111000,
	240'b101101101111111111100001011101101110001111111111111111111111111111111111111111111111111111111111111111111111111111110110110001110111111001010011010100110101010001010001010101110101101101010011010100100101001101100000111000101111111010111000,
	240'b101101101111111111100001101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110110001011000000101000101010101010101000101010001010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111101100111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010111000101010000010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111110011111110101111111111111111111111111111111111111111111111111111111111111111111111111111010011101001111010011111010011111111111111111110011101111101010100000101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111110100111110011111111111111111111111111111111111111111111111111111111111100010100111110111001101100001011000010111001110011111111000101111111111101100011111000101000001010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111110010111110011111111111111111111111111111111111111111111111111100001001100110010011110100111001001101010011010100111001001111011001101100000111111111111001010110110101010001010101010101001101100000111000101111111010111000,
	240'b101101101111111111101110111100101111111111111111111111111111111111111111110001110101101001010001010110000111010010010000100100000111010001010100010011110101101011000100111111111100110101011011010100110101001101100000111000101111111010111000,
	240'b101101101111111111101000111000001111111111111111111111111111111111101010011010110101000101010010011100101110101011111111111111111111001010110100010111100100111101101001111010001111111110100010010100010101001101100000111000101111111010111000,
	240'b101101101111111111100001110010011111111111111111111111111111111110101001010100000101001101010010010101011010000111111101111111111111111111111111101111100101011101001110101001001111111111101111011100000101000001100000111000101111111010111000,
	240'b101101101111111111011111101001111111111111111111111111111111011101110110010011100111100101110100010100000101010010101101111111111111111111111111111111011000100001001101011100101111010111111111101110010101000101100000111000101111111010111000,
	240'b101101101111111111100000100000111111011111111111111111111110001001011110010100001011111011100001011010100100111101011000101110111111111111111111111111111100000001010000010110111110000011111111111100010110110101011101111000101111111010111000,
	240'b101101101111111111100011011001111101100011111111111111111101010101010101010101011101011111111111110100010110001001001111010111011100100011111111111111111101100001011000010101101101000011111111111111111010011001011011111000101111111010111000,
	240'b101101101111111111100100010111001010010011111111111111111101010001010100010101011101100011111111111111111100010101011100010011110110010011010101111111111101100001011001010101101100111111111111111111111101100101100110111000001111111010111000,
	240'b101101101111111111100100010111100110110011110001111111111110000001011101010100011011111011111111111111111111111110111000010101110100111101101100111001001100011001010001010110101101111011111111111111111111011110000100110111101111111010111000,
	240'b101101101111111111100100011000000101000110110111111111111111010101110011010011001000100111111101111111111111111111111110101010100101001101001111011110010111111101001111011011111111001111111111111111111111111110101000110111001111111010111000,
	240'b101101101111111111100100011000010101000001101111111011111111111110100100010011100101100011000011111111111111111111111111111111001001111101010101010100100101001101010000101000001111111111111111111111111111111111001010111000001111110110111000,
	240'b101101101111111111100100011000010101001101010001101000101111111111100110011001110100111101100001101111101111100011111111111111111111000001110110010100100101000101100101111001001111111111111111111111111111111111100011111001001111110110111000,
	240'b101101101111111111100100011000010101001101010011010111001101000111111111110000000101011101010000010101110111110010011010100110110111110101011010010100010101011010111011111111111111111111111111111111111111111111110000111010111111110010111000,
	240'b101101101111111111100100011000010101001101010101010100010110111111100110111111111011100101100000010011100100111001001111010011110100111001001111010111111011011011111110111111111111111111111111111111111111111111110100111100011111110010111000,
	240'b101101101111111111100100011000010101001101010101010101010101000010000000111011101111111111011001100100110110100101011101010111010110011110010001110110001111111111111111111111111111111111111111111111111111111111110110111101001111110010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010000100000111110110011111111111111111110111011011100110110111110110111111110111111111111111111111111111111111111111111111111111111111111111111110110111100111111101110111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010100010111011111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111010111111110010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010001010100010101010101000001100101101110011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101110111111111111010111000,
	240'b101101101111111111100100011000010101001101010011010100010101011101010011010100010101010101010010010101011000010011001101111110011111111111111111111111111111111111111111111111111111111111111111111111111110100101111100110111101111111010111000,
	240'b101101101111111111100100011000010101000001100011101010001100111011000100100001000101010001010101010101000101000101011001011111111011100011100010111110001111111111111111111111111111111111111111111001001000000001011100111000101111111010111000,
	240'b101101101111111111100100010111110110000011010011111100111100001111010101111101011001010101010001010101010101010101010100010100010101001101100000011111001001001010101000101100111011010010011001011010000101000001100000111000101111111010111000,
	240'b101101101111111111100100010111011010001111111111111010110111000001010001101011011110101001101000010100110101010101010101010101010101010101010011010100010101000001010001010100100101001001010000010100100101001101100000111000101111111010111000,
	240'b101101101111111111100011011000111101010110111000110100011101111101100100010111111110100110001110010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111100011011001111101111110010101011001001110001011010001011001011110000010011000010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111100100011000001100101011000001010011000111000011100101110101101110110110000000010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111100100010111001000011111110110101001000110010110100010111111111101001001011011010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101011111111111011101101011001000101001010100011111100101110111111110000110101100111000001010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100100111010011111111010101101,
	240'b100111111111000111111101100101110100110101001110011011101001000010000100010110100100110101010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111010010100111111011111011010011011,
	240'b110001011101010111111111111100101010100010001000100001101000010010000101100010001000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010011010011111110000111111111101011011000101,
	240'b111111001100001111100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001100001111111100,
	240'b111101101110101110111111110110001110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011011000101110101110100111110110,
	240'b111011101111001111110011101001101000110010101001101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010101000110110011100111001001111000111101110,
	240'b111111111111111111100111101000001001110010110111101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110001001110110100110111100111111111111111111,
	240'b111111111111011010111011110011011110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011010000110000011111011011111111,
	240'b111111011100010111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100010011111101,
	240'b110010101101001011111111111101011011010110010101100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010011100100001000111110010001100101011011010011110100111111111101001111001010,
	240'b100111111111000011111110100111100100111101010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100010100111001010110011110001000010001100111010011010100111010011011111111101111010110011011,
	240'b101011101111111011101110011001100101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110100011001011111100111111001011101111100111000101000101100100111010111111111010101100,
	240'b101101101111111111100100011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101111100011111111111101010010111000110101111111101101000010001011011111000101111111010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011110011110111111011110110111110110101001001110110001001100100101011111111000011111111010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100101011101111101101110110101111101110001011111100100111101111001101001111000001111111010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100011001110100001100000011001111110001111001010101011111101100001100110111000001111111010111000,
	240'b101101101111111111100100011000010101001101010011010100000101000001010000010011110101000001010010010101000101010101010101010101010101010101010010011010001110110010101000010011110111000111101000111111101010110101011100111000011111111010111000,
	240'b101101101111111111100100011000010100111101100000100010111010010010100011100110011000100001110001010110110101000101010001010101000101010101010101010100101001101111110111110010111011001011110000110111100110010101011110111000101111111010111000,
	240'b101101101111111111100100010111010111011011011000111111101111111111111111111111111111110111110010110110001010111001111010010101100101000101010101010101000101010110001110110011111101110010110101011010100101000001100000111000101111111010111000,
	240'b101101101111111111100001011101101110001111111111111111111111111111111111111111111111111111111111111111111111111111110110110001110111111001010011010100110101010001010001010101110101101101010011010100100101001101100000111000101111111010111000,
	240'b101101101111111111100001101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110110001011000000101000101010101010101000101010001010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111101100111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010111000101010000010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111110011111110101111111111111111111111111111111111111111111111111111111111111111111111111111010011101001111010011111010011111111111111111110011101111101010100000101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111110100111110011111111111111111111111111111111111111111111111111111111111100010100111110111001101100001011000010111001110011111111000101111111111101100011111000101000001010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111110010111110011111111111111111111111111111111111111111111111111100001001100110010011110100111001001101010011010100111001001111011001101100000111111111111001010110110101010001010101010101001101100000111000101111111010111000,
	240'b101101101111111111101110111100101111111111111111111111111111111111111111110001110101101001010001010110000111010010010000100100000111010001010100010011110101101011000100111111111100110101011011010100110101001101100000111000101111111010111000,
	240'b101101101111111111101000111000001111111111111111111111111111111111101010011010110101000101010010011100101110101011111111111111111111001010110100010111100100111101101001111010001111111110100010010100010101001101100000111000101111111010111000,
	240'b101101101111111111100001110010011111111111111111111111111111111110101001010100000101001101010010010101011010000111111101111111111111111111111111101111100101011101001110101001001111111111101111011100000101000001100000111000101111111010111000,
	240'b101101101111111111011111101001111111111111111111111111111111011101110110010011100111100101110100010100000101010010101101111111111111111111111111111111011000100001001101011100101111010111111111101110010101000101100000111000101111111010111000,
	240'b101101101111111111100000100000111111011111111111111111111110001001011110010100001011111011100001011010100100111101011000101110111111111111111111111111111100000001010000010110111110000011111111111100010110110101011101111000101111111010111000,
	240'b101101101111111111100011011001111101100011111111111111111101010101010101010101011101011111111111110100010110001001001111010111011100100011111111111111111101100001011000010101101101000011111111111111111010011001011011111000101111111010111000,
	240'b101101101111111111100100010111001010010011111111111111111101010001010100010101011101100011111111111111111100010101011100010011110110010011010101111111111101100001011001010101101100111111111111111111111101100101100110111000001111111010111000,
	240'b101101101111111111100100010111100110110011110001111111111110000001011101010100011011111011111111111111111111111110111000010101110100111101101100111001001100011001010001010110101101111011111111111111111111011110000100110111101111111010111000,
	240'b101101101111111111100100011000000101000110110111111111111111010101110011010011001000100111111101111111111111111111111110101010100101001101001111011110010111111101001111011011111111001111111111111111111111111110101000110111001111111010111000,
	240'b101101101111111111100100011000010101000001101111111011111111111110100100010011100101100011000011111111111111111111111111111111001001111101010101010100100101001101010000101000001111111111111111111111111111111111001010111000001111110110111000,
	240'b101101101111111111100100011000010101001101010001101000101111111111100110011001110100111101100001101111101111100011111111111111111111000001110110010100100101000101100101111001001111111111111111111111111111111111100011111001001111110110111000,
	240'b101101101111111111100100011000010101001101010011010111001101000111111111110000000101011101010000010101110111110010011010100110110111110101011010010100010101011010111011111111111111111111111111111111111111111111110000111010111111110010111000,
	240'b101101101111111111100100011000010101001101010101010100010110111111100110111111111011100101100000010011100100111001001111010011110100111001001111010111111011011011111110111111111111111111111111111111111111111111110100111100011111110010111000,
	240'b101101101111111111100100011000010101001101010101010101010101000010000000111011101111111111011001100100110110100101011101010111010110011110010001110110001111111111111111111111111111111111111111111111111111111111110110111101001111110010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010000100000111110110011111111111111111110111011011100110110111110110111111110111111111111111111111111111111111111111111111111111111111111111111110110111100111111101110111000,
	240'b101101101111111111100100011000010101001101010101010101010101010101010101010100010111011111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111010111111110010111000,
	240'b101101101111111111100100011000010101001101010101010101010101010001010100010101010101000001100101101110011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101110111111111111010111000,
	240'b101101101111111111100100011000010101001101010011010100010101011101010011010100010101010101010010010101011000010011001101111110011111111111111111111111111111111111111111111111111111111111111111111111111110100101111100110111101111111010111000,
	240'b101101101111111111100100011000010101000001100011101010001100111011000100100001000101010001010101010101000101000101011001011111111011100011100010111110001111111111111111111111111111111111111111111001001000000001011100111000101111111010111000,
	240'b101101101111111111100100010111110110000011010011111100111100001111010101111101011001010101010001010101010101010101010100010100010101001101100000011111001001001010101000101100111011010010011001011010000101000001100000111000101111111010111000,
	240'b101101101111111111100100010111011010001111111111111010110111000001010001101011011110101001101000010100110101010101010101010101010101010101010011010100010101000001010001010100100101001001010000010100100101001101100000111000101111111010111000,
	240'b101101101111111111100011011000111101010110111000110100011101111101100100010111111110100110001110010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111100011011001111101111110010101011001001110001011010001011001011110000010011000010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111100100011000001100101011000001010011000111000011100101110101101110110110000000010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101101101111111111100100010111001000011111110110101001000110010110100010111111111101001001011011010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111010111000,
	240'b101011111111111011101101011001000101001010100011111100101110111111110000110101100111000001010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100100111010011111111010101101,
	240'b100111111111000111111101100101110100110101001110011011101001000010000100010110100100110101010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111010010100111111011111011010011011,
	240'b110001011101010111111111111100101010100010001000100001101000010010000101100010001000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010011010011111110000111111111101011011000101,
	240'b111111001100001111100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001100001111111100,
	240'b111101101110101110111111110110001110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011011000101110101110100111110110,
	240'b111011101111001111110011101001101000110010101001101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010101000110110011100111001001111000111101110,
	240'b111111111111111111100111101000001001110010110111101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110001001110110100110111100111111111111111111,
	240'b111111111111011010111011110011011110110011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110110011010000110000011111011011111111,
	240'b111111011100010111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100010011111101,
	240'b110010101101001011111111111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111111101001111001010,
	240'b100111111110111111111111111111101111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111101111111011111101111111011111110111111110111111111111010010011011,
	240'b101011101111110011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111110111111111111111111111111111111101111110111111101111111111111110010101100,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111011111111111111101111110111111110111111111111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111111111111111111110111111101111111101111111011111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111101111111111111111111111101111111101111111111111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111101111111011111111111111110111111101111111111111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111110111111011111110111111111111111111111111011111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111101111111011111110111111101111111011111101111111011111110111111101111111011111110111111101111111011111111011111111111111101111111011111111111111111111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111011111101111111011111110111111101111111011111110111111110111111101111111011111110111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111101111111011111110111111110111111111111111111111111111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111011111101111111011111110111111101111111011111110111111101111111011111111011111111111111111111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111101111110111111101111111011111110111111110111111101111110111111101111111011111110111111110111111111111111011111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111011111110111111101111111011111111111111111111111111111111111111110111111011111110111111101111111111111111111111110111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111101111111111111111111111111111111111111110111111011111110111111101111111011111111011111111111111111111111111111111111111101111110111111101111111101111111111111111111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111101111111111111111111111111111111111111101111111011111110111111101111111011111110111111110111111111111111111111111111111111111111011111101111111011111111111111111111111101111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111111111111111111111111111111111101111111011111111011111111111111011111110111111101111111101111111111111111111111111111111011111101111111011111111111111111111111111111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111111111111111111111111111111111101111111011111111011111111111111101111110111111101111111011111111011111111111111111111111111111101111111011111111011111111111111111111111011111101111111111111101010111000,
	240'b101101101111111011111111111111011111111011111111111111111111111111111101111111011111111011111111111111111111111011111101111111011111110111111111111111111111111011111101111111011111111011111111111111111111111011111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111111111111111111111111111101111111011111111011111111111111111111111111111110111111011111110111111101111111111111111011111101111111011111111111111111111111111111111111111110111111111111101010111000,
	240'b101101101111111011111111111111011111110111111110111111111111111111111101111111011111111011111111111111111111111111111111111111101111110111111101111111011111110111111101111111011111111111111111111111111111111111111110111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111111111111111111110111111011111110111111110111111111111111111111111111111111111111011111101111111011111110111111101111111101111111111111111111111111111111111111110111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111101111111111111111111111011111110111111101111111101111111111111111111111111111111111111101111111011111110111111101111111111111111111111111111111111111111111111111111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111111011111111111111101111110111111101111111011111111011111110111111101111110111111101111111011111110111111110111111111111111111111111111111111111111111111111111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111111111111111111111011111101111111011111110111111101111111011111110111111101111111011111111011111111111111111111111111111111111111111111111111111111111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111111111111111111110111111101111110111111101111111011111110111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111101111111101111111111111110111111011111110111111101111111011111110111111101111111011111111011111111111111111111111111111111111111111111111111111111111111111111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111110111111111111111111111111011111111111111111111111011111101111111011111110111111101111111011111110111111101111111101111111011111110111111101111111011111110111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111011111111111111111111110111111101111111101111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111111111110111111111111111111111101111111011111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111111111110111111011111111111111111111111011111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111111111110111111011111110111111111111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101101101111111011111111111111011111111011111111111111101111110111111110111111111111111011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101010111000,
	240'b101011111111110111111111111111011111110111111110111111111111111111111111111111101111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110101101,
	240'b100111111111000111111111111111101111110111111101111111011111111011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111010110011011,
	240'b110001011101010111111111111111111111111011111110111111101111110111111101111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111111101011011000101,
	240'b111111001100001111100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001100001111111100,
	240'b111101101110101110111111110110001110111011101110111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101110111011011000101110101110100111110110,
	240'b111011101111001111110011101001101000110010101001101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010101000110110011100111001001111000111101110,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule