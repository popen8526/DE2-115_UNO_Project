module blue_draw_two(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111111111111111111100100101000011001101110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001001001101010101100111100111111111111111111,
	240'b111111111110101110111001111000011111110011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111101111011110101111011110111111111111,
	240'b111101101011111111110010111111111111111111110111111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101111111111111111111111011011100000111111000,
	240'b101111001101111011111111111001011001001101111001011110000111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011101100111010001110100011101110111100101111000011110011001100011101010111111111101100010111010,
	240'b101000101111100111111010100001010100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111011010111010000010010000010110000101000001010001010100010100110110010000111111011111001110100001,
	240'b101011101111111111100100010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101111111001101110111011110111101110010101011001010100010101000101001001100110111011011111111010110000,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010101111110111110110100110010000111110000111010001010001010110000101010101100011111001111111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010111110110010100100110101011010101000000110100101010011101110011000000001011110111001111111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110001101111100111001001101010001010011010101110110011101111100111100011010001010111001011111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010001010100010101010101010101010101010101010101010101010101010101010101010101010011101000101111010110101100010110000110011011100000111111011111001110110110111000111111111010110100,
	240'b101100011111111111011110010111100101001101010010010100000101001101010011010100000101000001010001010100100101010001010101010101010101010001110011011100001001011011110010110010110110010001101000111001011010000001101001111001111111111010110100,
	240'b101100011111111111011110010111010101000001110001101001111011111110111110101101001010000010000100011001100101010001010000010100110101000011000000111011001100010111101011111111111000000001010000100001100110100001100001111001111111111010110100,
	240'b101100011111111111011110010110111000111011101100111111111111111111111111111111111111111111111100111010011100010010001101010111010100110110011001110010101100101011000111110000110111000101010010010100010101000101100100111001111111111010110100,
	240'b101100011111111111011010100001001111001011111111111111111111111111111111111111111111111111111111111111111111111111111110110110011000111001010110010100010101010001010100010101000101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011101110011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000010011010010101000001010100010101000101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111101010111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010111110101010001010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111011110010111110001111111111111111111111111110111111001000110001111100100011001000110010001100110111101100111111111111111111111111111111111110111110001000010100010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111011110001111101111111111111111111111111111100000111011110111100011110011111100110111010101110101011000011111100101111111111111111111111111111111111110001100001000101000001010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111101110111101101111111111111111111111111101000011101110101011110111000001110010011101011011101111100001110101111111111111111111111111111111111111111111111010100111001001010001010101010101001101100100111001111111111010110100,
	240'b101100011111111111101001111100101111111111111111111111111110000111011000100010100100110001010001010011110110000111010110110011101111111111111111111111111111111111111111111111111101001101011101010100110101001101100100111001111111111010110100,
	240'b101100011111111111100011111000111111111111111111111111111111001111001110101011100101000101010101010101010101001011000001101111001100100111001111110101111111010111111111111111111111111110100111010100010101001101100100111001111111111010110100,
	240'b101100011111111111011100110010101111111111111111111111111111110111001011110011010101100001010100010101010100111110011100110011101100111111101001110111101100010111111010111111111111111111110001011100010100111101100100111001111111111010110100,
	240'b101100011111111111011000101010001111111111111111111111111111111111010010110110010110110101010010010101010101000101111010110101110111101010000111110101101101010111100101111111111111111111111111101110100101000101100011111001111111111010110100,
	240'b101100011111111111011010100000111111100011111111111111111111111111100011110101111000110001010000010101010101001101011111110110010110110001001001011101101101110011010110111111111111111111111111111100010110110101100001111001111111111010110100,
	240'b101100011111111111011100011001011101101011111111111111111111111111110010110011111011000101010000010101010101010101010010110000011001011101001100010110111101000011001011111111101111111111111111111111111010010101011111111001111111111010110100,
	240'b101100011111111111011110010110011010011011111111111111111111111111111110110010111100110101011000010101000101010101010000100111001011101101001110010100011011011011001101111101011111111111111111111111111101011001101001111001101111111010110100,
	240'b101100011111111111011110010110110110110111110001111111111111111111111111110100111101110001110100010011000100111101001011011110101101110001011000010011111001001011010110111001101111111111111111111111111111010110000101111000111111111010110100,
	240'b101100011111111111011110010111010101000110110111111111111111111111111111111000101101011011011100100111001001100110011000110000011111101001101111010011010111000111011001110101001111111111111111111111111111111110101000111000011111111010110100,
	240'b101100011111111111011110010111100101000001101110111011101111111111111111111110111100011111011101111010001110011011100101111001011100111101100011010100010101101011001111110010111111111011111111111111111111111111001001111001001111111010110100,
	240'b101100011111111111011110010111100101001101010001101000011111111111111111111111111111100111011011110101101101000110101110101001010100111101010001010101010101000110110011110011011111010111111111111111111111111111100001111010011111110110110100,
	240'b101100011111111111011110010111100101001101010011010110111100111111111111111111111111111111111111111111111111111111001111110101110101111101001110010100000100101010010011110101111110001111111111111111111111111111110010111011101111110110110100,
	240'b101100011111111111011110010111100101001101010101010100010110110111100101111111111111111111111111111111111111111111010100111000111100010110001110100011101000110111001000111011011101000011111111111111111111111111110110111100011111110010110100,
	240'b101100011111111111011110010111100101001101010101010101010101000001111110111011001111111111111111111111111111111111110010110000101110010011100011111000101110001111100110110100011100100111111111111111111111111111110111111101001111110010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010000100000011110101011111111111111111111111111111111111100001101000011001111110100001101000011001110110100011111011111111111111111111111111111110111111100111111110010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010100010111010011011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111011011111110110110100,
	240'b101100011111111111011110010111100101001101010101010101010101010001010011010100110100111101100001101101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111001001111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101100001011101010111010101111001011011010110000111111111001001111101111111111111111111111111111111111111111111111111111111111111111111111111111110000001110111111001001111111010110100,
	240'b101100011111111111011110010111100101000101010010010100010111111111011000110110011101110011011101100111000100110001010111011110111011001111011110111101011111111111111111111111111111111111111111110110100111010101100000111001111111111010110100,
	240'b101100011111111111011110010110100111011010010000010011101000101111111111110111101011000011100010101011100101000001010100010100010101001001011110011101101000110010100001101010111010110010001111011000100100111101100100111001111111111010110100,
	240'b101100011111111111011110011011011011011011100010011100000110010011000000111100011001110101100110011000100101010001010101010101010101010101010011010100010101000001010001010100010101000101010000010100110101001101100100111001111111111010110100,
	240'b101100011111111111011100101111111111100111111101110111110110000101010101101000101111010010101101010101010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011101011111001100010011101000100001100101100101010000010100001000101011110011100010110101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011110010110001000001010100100010011100111100010110011010110010100111111010010101100110100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011110010111100101001001010011010100010111100111111000100101100111110111101101100111000101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101011011111111111100111011000010101001001010101010101000101011010110101111101101111010111010001011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111011111111110110101111,
	240'b101000001111011011111100100100010100111001010000010100000100111101010100100000001000100001011100010011100101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111110011100111111101111000010011111,
	240'b110001101101011111111111111100001010011110001011100011001000110010001011100001111000011110001010100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100010111010110011110100111111111101001011000101,
	240'b111111001100000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001100010011111101,
	240'b111101101110100010111110110110101111000011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101011110111111010101101110111110101111110101,
	240'b111011101111001011101111101000101000110110101010101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101010011000110010100001111001101111000111101110,
	240'b111111111111111111100100101000011001101110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001001001101010101100111100111111111111111111,
	240'b111111111110101110111001111000011111110011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111101111011110101111011110111111111111,
	240'b111101101011111111110010111111111111111111110111111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101111111111111111111111011011100000111111000,
	240'b101111001101111011111111111001011001001101111001011110000111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011101100111010001110100011101110111100101111000011110011001100011101010111111111101100010111010,
	240'b101000101111100111111010100001010100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111011010111010000010010000010110000101000001010001010100010100110110010000111111011111001110100001,
	240'b101011101111111111100100010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101111111001101110111011110111101110010101011001010100010101000101001001100110111011011111111010110000,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010101111110111110110100110010000111110000111010001010001010110000101010101100011111001111111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010111110110010100100110101011010101000000110100101010011101110011000000001011110111001111111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110001101111100111001001101010001010011010101110110011101111100111100011010001010111001011111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010001010100010101010101010101010101010101010101010101010101010101010101010101010011101000101111010110101100010110000110011011100000111111011111001110110110111000111111111010110100,
	240'b101100011111111111011110010111100101001101010010010100000101001101010011010100000101000001010001010100100101010001010101010101010101010001110011011100001001011011110010110010110110010001101000111001011010000001101001111001111111111010110100,
	240'b101100011111111111011110010111010101000001110001101001111011111110111110101101001010000010000100011001100101010001010000010100110101000011000000111011001100010111101011111111111000000001010000100001100110100001100001111001111111111010110100,
	240'b101100011111111111011110010110111000111011101100111111111111111111111111111111111111111111111100111010011100010010001101010111010100110110011001110010101100101011000111110000110111000101010010010100010101000101100100111001111111111010110100,
	240'b101100011111111111011010100001001111001011111111111111111111111111111111111111111111111111111111111111111111111111111110110110011000111001010110010100010101010001010100010101000101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011101110011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000010011010010101000001010100010101000101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111101010111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010111110101010001010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111011110010111110001111111111111111111111111110111111001000110001111100100011001000110010001100110111101100111111111111111111111111111111111110111110001000010100010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111011110001111101111111111111111111111111111100000111011110111100011110011111100110111010101110101011000011111100101111111111111111111111111111111111110001100001000101000001010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111101110111101101111111111111111111111111101000011101110101011110111000001110010011101011011101111100001110101111111111111111111111111111111111111111111111010100111001001010001010101010101001101100100111001111111111010110100,
	240'b101100011111111111101001111100101111111111111111111111111110000111011000100010100100110001010001010011110110000111010110110011101111111111111111111111111111111111111111111111111101001101011101010100110101001101100100111001111111111010110100,
	240'b101100011111111111100011111000111111111111111111111111111111001111001110101011100101000101010101010101010101001011000001101111001100100111001111110101111111010111111111111111111111111110100111010100010101001101100100111001111111111010110100,
	240'b101100011111111111011100110010101111111111111111111111111111110111001011110011010101100001010100010101010100111110011100110011101100111111101001110111101100010111111010111111111111111111110001011100010100111101100100111001111111111010110100,
	240'b101100011111111111011000101010001111111111111111111111111111111111010010110110010110110101010010010101010101000101111010110101110111101010000111110101101101010111100101111111111111111111111111101110100101000101100011111001111111111010110100,
	240'b101100011111111111011010100000111111100011111111111111111111111111100011110101111000110001010000010101010101001101011111110110010110110001001001011101101101110011010110111111111111111111111111111100010110110101100001111001111111111010110100,
	240'b101100011111111111011100011001011101101011111111111111111111111111110010110011111011000101010000010101010101010101010010110000011001011101001100010110111101000011001011111111101111111111111111111111111010010101011111111001111111111010110100,
	240'b101100011111111111011110010110011010011011111111111111111111111111111110110010111100110101011000010101000101010101010000100111001011101101001110010100011011011011001101111101011111111111111111111111111101011001101001111001101111111010110100,
	240'b101100011111111111011110010110110110110111110001111111111111111111111111110100111101110001110100010011000100111101001011011110101101110001011000010011111001001011010110111001101111111111111111111111111111010110000101111000111111111010110100,
	240'b101100011111111111011110010111010101000110110111111111111111111111111111111000101101011011011100100111001001100110011000110000011111101001101111010011010111000111011001110101001111111111111111111111111111111110101000111000011111111010110100,
	240'b101100011111111111011110010111100101000001101110111011101111111111111111111110111100011111011101111010001110011011100101111001011100111101100011010100010101101011001111110010111111111011111111111111111111111111001001111001001111111010110100,
	240'b101100011111111111011110010111100101001101010001101000011111111111111111111111111111100111011011110101101101000110101110101001010100111101010001010101010101000110110011110011011111010111111111111111111111111111100001111010011111110110110100,
	240'b101100011111111111011110010111100101001101010011010110111100111111111111111111111111111111111111111111111111111111001111110101110101111101001110010100000100101010010011110101111110001111111111111111111111111111110010111011101111110110110100,
	240'b101100011111111111011110010111100101001101010101010100010110110111100101111111111111111111111111111111111111111111010100111000111100010110001110100011101000110111001000111011011101000011111111111111111111111111110110111100011111110010110100,
	240'b101100011111111111011110010111100101001101010101010101010101000001111110111011001111111111111111111111111111111111110010110000101110010011100011111000101110001111100110110100011100100111111111111111111111111111110111111101001111110010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010000100000011110101011111111111111111111111111111111111100001101000011001111110100001101000011001110110100011111011111111111111111111111111111110111111100111111110010110100,
	240'b101100011111111111011110010111100101001101010101010101010101010101010101010100010111010011011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111011011111110110110100,
	240'b101100011111111111011110010111100101001101010101010101010101010001010011010100110100111101100001101101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111001001111111010110100,
	240'b101100011111111111011110010111100101001101010101010101010101100001011101010111010101111001011011010110000111111111001001111101111111111111111111111111111111111111111111111111111111111111111111111111111110000001110111111001001111111010110100,
	240'b101100011111111111011110010111100101000101010010010100010111111111011000110110011101110011011101100111000100110001010111011110111011001111011110111101011111111111111111111111111111111111111111110110100111010101100000111001111111111010110100,
	240'b101100011111111111011110010110100111011010010000010011101000101111111111110111101011000011100010101011100101000001010100010100010101001001011110011101101000110010100001101010111010110010001111011000100100111101100100111001111111111010110100,
	240'b101100011111111111011110011011011011011011100010011100000110010011000000111100011001110101100110011000100101010001010101010101010101010101010011010100010101000001010001010100010101000101010000010100110101001101100100111001111111111010110100,
	240'b101100011111111111011100101111111111100111111101110111110110000101010101101000101111010010101101010101010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011101011111001100010011101000100001100101100101010000010100001000101011110011100010110101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011110010110001000001010100100010011100111100010110011010110010100111111010010101100110100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101100011111111111011110010111100101001001010011010100010111100111111000100101100111110111101101100111000101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111001111111111010110100,
	240'b101011011111111111100111011000010101001001010101010101000101011010110101111101101111010111010001011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111011111111110110101111,
	240'b101000001111011011111100100100010100111001010000010100000100111101010100100000001000100001011100010011100101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111110011100111111101111000010011111,
	240'b110001101101011111111111111100001010011110001011100011001000110010001011100001111000011110001010100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100010111010110011110100111111111101001011000101,
	240'b111111001100000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001100010011111101,
	240'b111101101110100010111110110110101111000011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101011110111111010101101110111110101111110101,
	240'b111011101111001011101111101000101000110110101010101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101010011000110010100001111001101111000111101110,
	240'b111111111111111111100100101000011001101110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001001001101010101100111100111111111111111111,
	240'b111111111110101110111001111000011111110011111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111011110101111011110111111111111,
	240'b111101101011111111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011100000111111000,
	240'b101111001101111011111111111111111111111011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111011111111111111111101100010111010,
	240'b101000101111100011111111111111101111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111011111110111111011111110111111101111111011111110111111110111111111111001010100001,
	240'b101011101111111011111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111111111111111111111101111110111111101111111011111110111111101111111111111101110110000,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111110111111111111110111111110111111111111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111110111111101111110111111101111111101111110111111101111111101111111011111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111110111111111111111011111101111111011111110111111110111111111111111011111110111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111110111111011111110111111111111111111111111111111110111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111011111111111111101111110111111101111111111111111011111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111101111111011111110111111101111111011111110111111011111110111111101111111011111110111111110111111111111111011111111111111111111110111111101111111101111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111111011111111111111111111111111111111111111111111111111111111111111111111111011111110111111011111110111111110111111101111111011111110111111101111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111111111111111111111111111111110111111001000110001111100011111000111110001101100110111101100111111111111111111111111111111111111111111111110111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111111111111111111111111111111100000111011110111100011111000011110000111100011110100011000011111100101111111111111111111111111111111111111111111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111111111111111111111111111111100111111101101111111111111111111111111111111111111111111100001110101111111111111111111111111111111111111111111111111111111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111111111111111111111111111111110000011011000111111111111110111111101111111011111111111110001110010111111111111111111111111111111111111111111111111111111111111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111111111111111111111111111111111001011001001111111111111110111111101111111011111110111111110101101111100100011001110110101111111010111111111111111111111111111111110111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111101111111111111111111111111111110111000111111110001111111011111101111111011111110111111111110010111101000111101000110110111100010111111010111111111111111111111111111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111101111111111111111111111111111111111010000111010101111111111111101111111011111110111111111111000011101101011111111111111111101001111100101111111111111111111111111111111101111110111111101111111111111101110110100,
	240'b101100011111110111111111111111101111111111111111111111111111111111100010110101111111111111111101111111011111110111111110111101001100011111111111111111111110010111010100111111111111111111111111111111111111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111111111111111111111111111111111110010110010101111111011111101111111011111110111111101111111001100011111110101111111111111011011000110111111101111111111111111111111111111111011111101111111111111101110110100,
	240'b101100011111110111111111111111011111111011111111111111111111111111111110110001101111100011111110111111011111110111111101111111111101000011101000111111111111111011001000111101011111111111111111111111111111111111111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111111111111111111111111111111110100011110100011111111111111011111110111111101111111111110010011010011111111111111111111010100111001011111111111111111111111111111111111111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111110111111111111111111111111111000101101010011111111111111111111111111111111111111111111010011001000111111011111111111100111110100101111111111111111111111111111111111111110111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111111111111111111111111110101100011111011010111001011110010111100011111001101101011011000010111111011111111011110111110001111111111011111111111111111111111111111110111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111101111111111111111111111111111100111011011110101101101000110101010110101011101011011110011111111101111110111111111110010001111010111111111111111111111111111111110111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111111011111111111111111111111111111111111111111111111111001011111101111111111111111110111111011111110111111111110101011110001111111111111111111111111111111111111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111111111111111111111111111111111111111111111111010100111000111111111111111111111111111111111111111111111010111101000011111111111111111111111111111111111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111111111111111111111111111111111111111110010110000101110000111100100111001001110010011100100110100011100100111111111111111111111111111111111111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111111111111111111111111111111111111111111100001101000011001111110011111100111111001110110100011111011111111111111111111111111111111111111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111111011111111111111111111111111111111111111101111110111111101111111011111111011111111111111111111111111111111111111111111111111111111111111111111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111110111111011111111011111111111111101111111011111111111111101111110111111101111111011111110111111101111111011111111011111110111111101111111011111110111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111111011111111111111011111110111111110111111111111111011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111101111111111111111111111111111110111111101111111101111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111111011111111111111101111110111111101111111011111110111111111111111101111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111111011111110111111011111110111111110111111011111110111111111111111101111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101100011111110111111111111111011111110111111101111111011111110111111111111111101111111011111111111111101111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110110100,
	240'b101011011111110111111111111111011111110111111101111111011111110111111110111111111111111111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111101110101111,
	240'b101000001111010111111111111111101111110111111101111111011111110111111101111111011111111011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111110111111111110111110011111,
	240'b110001101101011111111111111111111111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111111111111101001011000101,
	240'b111111001100000111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001100010011111101,
	240'b111101101110100010111110110110101110111111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011110111111010101101110111110101111110101,
	240'b111011101111001011101111101000101000110110101010101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101010011000110010100001111001101111000111101110,
};
assign data = picture[addr];
endmodule