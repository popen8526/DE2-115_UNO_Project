module green_two(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111100111111111111101011101010001010010110101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101010001110100100111000111111001111110010,
	240'b111100111111011011000110110010101110010011110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011110001011000110101111101110100111110010,
	240'b111100011100001011100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011110111110001,
	240'b110001001101001111111111111101101011101010100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011001111010011100100111111011111011111000111111111100111011000101,
	240'b101000001111011011111101100110100101000001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011010110001001111000010111110100111010100010111111101111000110011110,
	240'b101010111111111111100110011000000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011111101110011111111011111000100111001001100010111011011111111110101101,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011001110101001100110001111101110101111100110001011111111000011111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100011111010101000111001000110100001011011011001100110111000011111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100011100110001011100010100010101011001100000111000101111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011100111110001011010010011011110100111001100000111000101111111110110100,
	240'b101100011111111111011001010111000101010001010011010100000100111101001111010100000101000101010010010101000101010101010101010101010101010101010101010101010101010101010111011000100110111111001111111001111000100101011111111000101111111110110100,
	240'b101100011111111111011001010111000101000001100000100010111010000110011110100101011000000001101010010110010101000001010010010101000101010101010101010101010101001101100011110111011011101110110100111110101110000101101001111000001111111110110011,
	240'b101100011111111111011001010110000111101011011010111111011111111111111111111111111111101011110000110100001010010001110001010101000101000101010101010101010101001101100010110100101110011111100101111000101100011001101000111000001111111110110011,
	240'b101100011111111111010110011101111110100011111111111111111111111111111111111111111111111111111111111111111111111111110001110000000111011001010010010100110101010101010110010110110101110001011100010111000101100101100000111000101111111110110011,
	240'b101100011111111111011000110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101001010111010101000101010101010101000101010001010100010101000101001001100000111000101111111110110011,
	240'b101100011111111111100110111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110110110101010001010101010101010101010101010101010101001101100000111000101111111110110011,
	240'b101100011111111111110000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111001111111000111111111111111111110010001111000010100000101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111110001111110001111111111111111111111111111111111111111111111111111111111111111111011001001110101101110011001000111000010100101111100011111111111100111011110000101000001010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111101110111101111111111111111111111111111111111111111111111111111111111111101000011110000100111101001110010011100100111001001111100000101111000011111111111000010110101101010010010101010101001101100000111000101111111110110100,
	240'b101100011111111111101000111101001111111111111111111111111111111111111111111111111111110110010011010011100101010001110111100101000111001001010010010011101010000111111111111111111100101001011010010101000101001101100000111000101111111110110100,
	240'b101100011111111111100010111001111111111111111111111111111111111111111111111111111110001001100000010100001000110111110010111111111110110110000010010011100110100011101100111111111111111110100000010100010101001101100000111000101111111110110100,
	240'b101100011111111111011010110100001111111111111111111111111111111111111111111111111100010101010001010110111101101011111111111111111111111111001101010100010101001011010010111111111111111111101101011011100101000001100000111000101111111110110100,
	240'b101100011111111111010100101011111111111111111111111111111111111111111111111111111011110101001110011000011110100011111111111111111111111111100110011111100111011111010100111111111111111111111111101101110101000101100000111000101111111110110011,
	240'b101100011111111111010101100010011111101111111111111111111111111111111111111111111100111001010101010101001100001111111111111111111111111111111101111101101111011011111100111111111111111111111111111100010110110101011101111000101111111110110011,
	240'b101100011111111111010111011001111110000111111111111111111111111111111111111111111111000001101101010011010111010011100100111111111111111111111111111111111111111111111111111111111111111111111111111111111010011001011011111000101111111110110011,
	240'b101100011111111111011001010110001011000011111111111111111111111111111111111111111111111110111100010101100100111101101110110100001111111111111111111111111111111111111111111111111111111111111111111111111101100101100110111000001111111110110011,
	240'b101100011111111111011001010110000111010011110110111111111111111111111111111111111111111111111101101101000101100001001110010111111011000011111010111111111111111111111111111111111111111111111111111111111111011110000100110111101111111110110011,
	240'b101100011111111111011001010110110101001111000000111111111111111111111111111111111111111111111111111111111011110101011111010011100101001110001100111001111111111111111111111111111111111111111111111111111111111110101001110111001111111110110100,
	240'b101100011111111111011001010111000101000001110101111100111111111111111111111111111111111111111111111111111111111111010010011100110100111101001111011011011100011111111101111111111111111111111111111111111111111111001010111000001111111110110100,
	240'b101100011111111111011001010111000101001101010010101010011111111111111111111111111101000110001001100110001111010111111111111011001000111001010110010100000101101111010100111111111111111111111111111111111111111111100011111001101111111110110100,
	240'b101100011111111111011001010111000101010001010011010111101101010111111111111111111011100001001001010101111001010110011111101000011001011101100000010100110101001111000111111111111111111111111111111111111111111111110011111011001111111110110100,
	240'b101100011111111111011001010111000101010001010101010100010111001011101001111111111011100101001101010100110100111101001110010011100100111101010011010100100101001011000111111111111111111111111111111111111111111111110111111100001111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101000010000001111100111100001101011011011000000110000001100000011000000110000001100000010111110110000011001100111111111111111111111111111111111111111111111000111100101111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010000100001011101111111100011111000011110000011100000111000001110000011100000111000001110000011110101111111111111111111111111111111111111111111111000111100101111111110110011,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010100000111100011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111010111111111110110011,
	240'b101100011111111111011001010111000101001101010100010101000101010001010100010101010101000101100011101100011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111111110110011,
	240'b101100011111111111011001010111010101101001011100010111000101110001011010010101010101010101010010010100110111101111000011111101011111111111111111111111111111111111111111111111111111111111111111111111111110001001110110110111111111111110110011,
	240'b101100011111111111011000011010001100100111011111111000011110001111001000010111010101001101010101010101000101000101010110011110001010111111011001111101011111110111111111111111111111111111111110110110100111011101011100111000101111111110110100,
	240'b101100011111111111010111011010101110110011110111101101001100011011011010010111100101001101010101010101010101010101010100010100010101000101011101011100011000100110011110101001111010100010001100011000000101000001100000111000101111111110110100,
	240'b101100011111111111011001010111001001011111101100110001000110101101100011010101100101010101010101010101010101010101010101010101010101010101010011010100100101000001010000010011110100111101010000010100110101001101100000111000101111111110110100,
	240'b101100011111111111011001010110110100111001111000110111111101110001101011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111011001010111000101010101010000011001001101100011000101010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111011000011001101011011101111011010001101001101011100011010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111011000010111111101100011001100011101101101000011001110010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110011,
	240'b101011001111111111100101010111000111111111101010111110011110011001111100010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100101111011001111111110101101,
	240'b100111111111011011111100100101100100110101100100011110110110001001001101010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101000010011111111111101111001010011101,
	240'b110000001101010111111111111101001011010010011001100110001001101010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001011100011110111111111111101000011000001,
	240'b111100001100000111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011101111110000,
	240'b111110011110110110111101110011001110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111000111111001,
	240'b111111001111001011011110100111111010001010110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100101010000110101001111100011111111111111101,
	240'b111100111111111111101011101010001010010110101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101010001110100100111000111111001111110010,
	240'b111100111111011011000110110010101110001111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011110001011000110101111101110100111110010,
	240'b111100011100001011100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011110111110001,
	240'b110001001101001111111111111110101101110111010000110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111011001101110011111101111011111100111111111100111011000101,
	240'b101000001111010111111110110011001010100010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001101011000010111011101011111010011111010001111111111111000110011110,
	240'b101010111111111111110010101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111111111001111111101111100001011100110110001111101101111111010101101,
	240'b101100011111111111101100101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101100111010011110011010111110111010111110010110101111111100001111111110110100,
	240'b101100011111111111101100101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110001111101001100011010100010110000101101101110110010111100001111111110110100,
	240'b101100011111111111101100101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101100111010001110010110101110101010001010101010101111111100001111111110110100,
	240'b101100011111111111101100101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111000111101001101101111010011010101111111100001111111110110100,
	240'b101100011111111111101100101011011010100110101001101010001010011110100111101001111010100010101001101010011010101010101010101010101010101010101010101010101010101010101011101100001011011111100111111100111100010010101111111100001111111110110100,
	240'b101100011111111111101100101011011010011110101111110001011101000011001111110010101100000010110100101011001010100010101000101010101010101010101010101010101010100110110001111011101101110111011001111111001111000010110100111100001111111110110011,
	240'b101100011111111111101100101010111011110111101100111111101111111111111111111111111111110111110111111001111101001010111000101010101010100010101010101010101010100110110000111010011111001111110010111100011110001010110011111100001111111110110011,
	240'b101100011111111111101011101110111111001111111111111111111111111111111111111111111111111111111111111111111111111111111000111000001011101010101000101010011010101010101010101011011010111010101110101011101010110010101111111100001111111110110011,
	240'b101100011111111111101100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011010100101011101010100010101010101010011010100110101001101010011010100010101111111100001111111110110011,
	240'b101100011111111111110011111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011011010101000101010101010101010101010101010101010100110101111111100001111111110110011,
	240'b101100011111111111111000111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111100111111100011111111111111111111000110111100101010001010101010101010101010101010100110101111111100001111111110110100,
	240'b101100011111111111111000111111001111111111111111111111111111111111111111111111111111111111111111111101101100111010110110101100101011100011010010111110001111111111110011101111001010100010101010101010101010100110101111111100001111111110110100,
	240'b101100011111111111110111111110111111111111111111111111111111111111111111111111111111111111110100101111001010011110100111101001101010011110100111110000011111011111111111111100001011010110101000101010101010100110101111111100001111111110110100,
	240'b101100011111111111110100111110101111111111111111111111111111111111111111111111111111111011001001101001111010100110111011110010011011100110101001101001111101000011111111111111111110010110101100101010011010100110101111111100001111111110110100,
	240'b101100011111111111110000111100111111111111111111111111111111111111111111111111111111000110101111101001111100011011111000111111111111011011000001101001111011001111110101111111111111111111001111101010001010100110101111111100001111111110110100,
	240'b101100011111111111101101111010001111111111111111111111111111111111111111111111111110001010101000101011011110110111111111111111111111111111100110101010001010100011101001111111111111111111110110101101101010011110101111111100001111111110110100,
	240'b101100011111111111101010110101111111111111111111111111111111111111111111111111111101111010100111101100001111001111111111111111111111111111110011101111111011101111101001111111111111111111111111110110111010100010101111111100001111111110110011,
	240'b101100011111111111101010110001001111110111111111111111111111111111111111111111111110011110101010101010101110000111111111111111111111111111111110111110111111101011111101111111111111111111111111111110001011011010101110111100001111111110110011,
	240'b101100011111111111101011101100111111000011111111111111111111111111111111111111111111100010110110101001101011101011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111101001010101101111100001111111110110011,
	240'b101100011111111111101100101010111101011111111111111111111111111111111111111111111111111111011101101010101010011110110111111010001111111111111111111111111111111111111111111111111111111111111111111111111110110010110011111100001111111110110011,
	240'b101100011111111111101100101010111011101011111010111111111111111111111111111111111111111111111110110110011010101110100110101011111101011111111100111111111111111111111111111111111111111111111111111111111111101111000001111011101111111110110011,
	240'b101100011111111111101100101011011010100111100000111111111111111111111111111111111111111111111111111111111101111010101111101001111010100111000101111100111111111111111111111111111111111111111111111111111111111111010100111011101111111110110100,
	240'b101100011111111111101100101011011010011110111010111110011111111111111111111111111111111111111111111111111111111111101000101110011010011110100111101101101110001111111110111111111111111111111111111111111111111111100101111011111111111110110100,
	240'b101100011111111111101100101011011010100110101000110101001111111111111111111111111110100011000100110010111111101011111111111101011100011010101011101010001010110111101001111111111111111111111111111111111111111111110001111100111111111110110100,
	240'b101100011111111111101100101011011010100110101001101011111110101011111111111111111101101110100100101010111100101011001111110100001100101110101111101010011010100111100010111111111111111111111111111111111111111111111001111101011111111110110100,
	240'b101100011111111111101100101011011010100110101010101010001011100011110100111111111101110010100110101010011010011110100110101001101010011110101001101010011010100111100011111111111111111111111111111111111111111111111011111101111111111010110100,
	240'b101100011111111111101100101011011010100110101010101010101010100011000000111110011110000110101101101100001011000010110000101100001011000010110000101100001011000011100101111111111111111111111111111111111111111111111011111110011111111010110100,
	240'b101100011111111111101100101011011010100110101010101010101010101010101000110000101110111111110001111100001111000011110000111100001111000011110000111100001111000011111010111111111111111111111111111111111111111111111100111110011111111010110011,
	240'b101100011111111111101100101011011010100110101010101010101010101010101010101010001011101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101011111111110110011,
	240'b101100011111111111101100101011011010100010101001101010011010100110101001101010101010100010110001110110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111011111111111110110011,
	240'b101100011111111111101100101011101010110010101101101011011010110110101101101010101010101010101001101010011011110111100001111110101111111111111111111111111111111111111111111111111111111111111111111111111111000110111010111011111111111110110011,
	240'b101100011111111111101011101101001110010011101110111100001111000111100011101011101010100110101010101010101010100010101011101111001101011111101100111110101111111011111111111111111111111111111110111011001011101110101101111100001111111110110100,
	240'b101100011111111111101011101101011111010111111011110110011110001011101100101011111010100110101010101010101010101010101010101010001010100010101110101110001100010011001110110100111101010011000101101011111010011110101111111100001111111110110100,
	240'b101100011111111111101100101011101100101111110110111000101011010110110001101010111010101010101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100110101111111100001111111110110100,
	240'b101100011111111111101100101011011010011110111100111011111110111010110101101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111111110110100,
	240'b101100011111111111101100101011011010101010101000101100011110101111100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111111110110100,
	240'b101100011111111111101011101100111101101110111101101000101100110011110001101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111111110110100,
	240'b101100011111111111101100101011111110110011100101101110101110011111100110101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111111110110011,
	240'b101011001111111111110010101011011011111111110100111111001111001110111110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101101111111110101101,
	240'b100111111111011011111110110010101010011010110001101111011011000110100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011111001111111111111111000110011101,
	240'b110000001101010111111111111110101101100111001100110010111100110011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011011101101111111011111111111101000011000001,
	240'b111100001100000111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011101111110000,
	240'b111110011110110110111101110011001110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111000111111001,
	240'b111111001111001011011110100111111010001010110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100101010000110101001111100011111111111111101,
	240'b111100111111111111101011101010001010010110101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101010001110100100111000111111001111110010,
	240'b111100111111011011000110110010101110010011110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011110001011000110101111101110100111110010,
	240'b111100011100001011100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011110111110001,
	240'b110001001101001111111111111101101011101010100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011001111010011100100111111011111011111000111111111100111011000101,
	240'b101000001111011011111101100110100101000001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011010110001001111000010111110100111010100010111111101111000110011110,
	240'b101010111111111111100110011000000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011111101110011111111011111000100111001001100010111011011111111110101101,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011001110101001100110001111101110101111100110001011111111000011111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100011111010101000111001000110100001011011011001100110111000011111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100011100110001011100010100010101011001100000111000101111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011100111110001011010010011011110100111001100000111000101111111110110100,
	240'b101100011111111111011001010111000101010001010011010100000100111101001111010100000101000101010010010101000101010101010101010101010101010101010101010101010101010101010111011000100110111111001111111001111000100101011111111000101111111110110100,
	240'b101100011111111111011001010111000101000001100000100010111010000110011110100101011000000001101010010110010101000001010010010101000101010101010101010101010101001101100011110111011011101110110100111110101110000101101001111000001111111110110011,
	240'b101100011111111111011001010110000111101011011010111111011111111111111111111111111111101011110000110100001010010001110001010101000101000101010101010101010101001101100010110100101110011111100101111000101100011001101000111000001111111110110011,
	240'b101100011111111111010110011101111110100011111111111111111111111111111111111111111111111111111111111111111111111111110001110000000111011001010010010100110101010101010110010110110101110001011100010111000101100101100000111000101111111110110011,
	240'b101100011111111111011000110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101001010111010101000101010101010101000101010001010100010101000101001001100000111000101111111110110011,
	240'b101100011111111111100110111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110110110101010001010101010101010101010101010101010101001101100000111000101111111110110011,
	240'b101100011111111111110000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111001111111000111111111111111111110010001111000010100000101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111110001111110001111111111111111111111111111111111111111111111111111111111111111111011001001110101101110011001000111000010100101111100011111111111100111011110000101000001010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111101110111101111111111111111111111111111111111111111111111111111111111111101000011110000100111101001110010011100100111001001111100000101111000011111111111000010110101101010010010101010101001101100000111000101111111110110100,
	240'b101100011111111111101000111101001111111111111111111111111111111111111111111111111111110110010011010011100101010001110111100101000111001001010010010011101010000111111111111111111100101001011010010101000101001101100000111000101111111110110100,
	240'b101100011111111111100010111001111111111111111111111111111111111111111111111111111110001001100000010100001000110111110010111111111110110110000010010011100110100011101100111111111111111110100000010100010101001101100000111000101111111110110100,
	240'b101100011111111111011010110100001111111111111111111111111111111111111111111111111100010101010001010110111101101011111111111111111111111111001101010100010101001011010010111111111111111111101101011011100101000001100000111000101111111110110100,
	240'b101100011111111111010100101011111111111111111111111111111111111111111111111111111011110101001110011000011110100011111111111111111111111111100110011111100111011111010100111111111111111111111111101101110101000101100000111000101111111110110011,
	240'b101100011111111111010101100010011111101111111111111111111111111111111111111111111100111001010101010101001100001111111111111111111111111111111101111101101111011011111100111111111111111111111111111100010110110101011101111000101111111110110011,
	240'b101100011111111111010111011001111110000111111111111111111111111111111111111111111111000001101101010011010111010011100100111111111111111111111111111111111111111111111111111111111111111111111111111111111010011001011011111000101111111110110011,
	240'b101100011111111111011001010110001011000011111111111111111111111111111111111111111111111110111100010101100100111101101110110100001111111111111111111111111111111111111111111111111111111111111111111111111101100101100110111000001111111110110011,
	240'b101100011111111111011001010110000111010011110110111111111111111111111111111111111111111111111101101101000101100001001110010111111011000011111010111111111111111111111111111111111111111111111111111111111111011110000100110111101111111110110011,
	240'b101100011111111111011001010110110101001111000000111111111111111111111111111111111111111111111111111111111011110101011111010011100101001110001100111001111111111111111111111111111111111111111111111111111111111110101001110111001111111110110100,
	240'b101100011111111111011001010111000101000001110101111100111111111111111111111111111111111111111111111111111111111111010010011100110100111101001111011011011100011111111101111111111111111111111111111111111111111111001010111000001111111110110100,
	240'b101100011111111111011001010111000101001101010010101010011111111111111111111111111101000110001001100110001111010111111111111011001000111001010110010100000101101111010100111111111111111111111111111111111111111111100011111001101111111110110100,
	240'b101100011111111111011001010111000101010001010011010111101101010111111111111111111011100001001001010101111001010110011111101000011001011101100000010100110101001111000111111111111111111111111111111111111111111111110011111011001111111110110100,
	240'b101100011111111111011001010111000101010001010101010100010111001011101001111111111011100101001101010100110100111101001110010011100100111101010011010100100101001011000111111111111111111111111111111111111111111111110111111100001111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101000010000001111100111100001101011011011000000110000001100000011000000110000001100000010111110110000011001100111111111111111111111111111111111111111111111000111100101111111110110100,
	240'b101100011111111111011001010111000101010001010101010101010101010101010000100001011101111111100011111000011110000011100000111000001110000011100000111000001110000011110101111111111111111111111111111111111111111111111000111100101111111110110011,
	240'b101100011111111111011001010111000101010001010101010101010101010101010101010100000111100011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111010111111111110110011,
	240'b101100011111111111011001010111000101001101010100010101000101010001010100010101010101000101100011101100011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111111110110011,
	240'b101100011111111111011001010111010101101001011100010111000101110001011010010101010101010101010010010100110111101111000011111101011111111111111111111111111111111111111111111111111111111111111111111111111110001001110110110111111111111110110011,
	240'b101100011111111111011000011010001100100111011111111000011110001111001000010111010101001101010101010101000101000101010110011110001010111111011001111101011111110111111111111111111111111111111110110110100111011101011100111000101111111110110100,
	240'b101100011111111111010111011010101110110011110111101101001100011011011010010111100101001101010101010101010101010101010100010100010101000101011101011100011000100110011110101001111010100010001100011000000101000001100000111000101111111110110100,
	240'b101100011111111111011001010111001001011111101100110001000110101101100011010101100101010101010101010101010101010101010101010101010101010101010011010100100101000001010000010011110100111101010000010100110101001101100000111000101111111110110100,
	240'b101100011111111111011001010110110100111001111000110111111101110001101011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111011001010111000101010101010000011001001101100011000101010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111011000011001101011011101111011010001101001101011100011010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110100,
	240'b101100011111111111011000010111111101100011001100011101101101000011001110010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111000101111111110110011,
	240'b101011001111111111100101010111000111111111101010111110011110011001111100010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100101111011001111111110101101,
	240'b100111111111011011111100100101100100110101100100011110110110001001001101010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101000010011111111111101111001010011101,
	240'b110000001101010111111111111101001011010010011001100110001001101010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001011100011110111111111111101000011000001,
	240'b111100001100000111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011101111110000,
	240'b111110011110110110111101110011001110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111000111111001,
	240'b111111001111001011011110100111111010001010110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100101010000110101001111100011111111111111101,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule