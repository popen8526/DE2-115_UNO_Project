module yellow_four(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110101111100011011110100101001001010110101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010001000110010110010111101011111101111111001,
	240'b111111111110100010111010110011001110000111101101111011101110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101110111010101101110011000101110100011111111111111110,
	240'b111110101011110011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101101010111111110,
	240'b110010111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100010111001010,
	240'b101000001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100110100000,
	240'b101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110101100,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101100001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110010,
	240'b101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110101111,
	240'b100111011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110100001,
	240'b101101111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101110110011,
	240'b111100001011110011111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100011111110101,
	240'b111111101101100110111100111010101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111101011011010101111111111010011111110,
	240'b111100011111111011100110101010011010001010101010101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101011101010111010101110101011101010001001111010110010111010111111001111110010,
	240'b111110101111100011011110100101001001010110101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010001000110010110010111101011111101111111001,
	240'b111111111110100010111010110011001110000111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101101110011000101110100011111111111111110,
	240'b111110101011110011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101101010111111110,
	240'b110010111101011111111111111110011101101011001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100110111001110110100001110011011111111111111011100010111001010,
	240'b101000001111101011111101110010001010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101010001011100110110001101001101010110011100001111111111101100110100000,
	240'b101001011111111111101110101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101110111100010101010101010011010111111111111111110101110101100,
	240'b101100001111111111101000101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111011101111110110101110101010011010111010111111001111010010110010,
	240'b101100001111111111101000101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101110111100110111101000110110011010011010111010111111001111010110110010,
	240'b101100001111111111101000101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110011101110111011000111111100101011000110111001111111001111010110110010,
	240'b101100001111111111101000101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110011101110111110110001111011111100110110111000111111001111010110110010,
	240'b101100001111111111101000101010111010101010101001101010001010011110101000101010001010100010101001101010101010101010101010101010101010101010101010101010101010100010110100111100011111110011101100111110111110010010111010111111001111010110110010,
	240'b101100011111111111101000101010111010100010101111110000101100110011001011110001101011101010110001101010011010100010101001101010101010101010101010101010101010100110110001111010011111101011011101110110111100100110111010111111001111010110110010,
	240'b101100011111111111101000101010011011110111101100111111101111111111111111111111111111110011110010111000011100100110110010101010001010100110101010101010101010101010100111110001111110001110101010101010011010011110111010111111001111010110110010,
	240'b101100011111111111100110101110101111010011111111111111111111111111111111111111111111111111111111111111111111111111110010110100111011001010101000101010101010101010101010101011011010111110101010101010101010100010111010111111001111010110110010,
	240'b101100011111111111101000111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011000110101010101010100110101010101010101010100110101010101010101010100010111010111111001111010110110010,
	240'b101100011111111111110001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110011010111010101000101010101010101010101010101010101010100010111010111111001111010110110010,
	240'b101100001111111111111000111111001111111111111111111111111111111111111111111111111111111111111111111111011111010111110101111110111111111111111111111111111110001110110000101010001010101010101010101010101010100010111010111111001111010110110010,
	240'b101100001111111111111001111111001111111111111111111111111111111111111111111111111111111111111111111110111100010010110010110100011111111111111111111111111111111111100101101100001010100110101010101010101010100010111010111111001111010110110010,
	240'b101100001111111111110111111110111111111111111111111111111111111111111111111111111111111111111111111111111101011010100101101100011111001111111111111111111111111111111111111000001010110010101001101010101010100010111010111111001111010110110010,
	240'b101100001111111111110100111110101111111111111111111111111111111111111111111111111111111111111111111111111111010010110010101001111101011111111111111111111111111111111111111111111101000110101000101010101010100010111010111111001111010110110010,
	240'b101100001111111111101110111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111001101101001101011100011111001111111111111111111111111111111111111100110111101101010001010100010111010111111001111010110110010,
	240'b101100001111111111101010111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101011011010100011100000111111111111111111111111111111111111111111100110101011001010011110111010111111001111010110110010,
	240'b101100011111111111100110110111011111111111111111111111111111111111111111111111111111111111110111110100111100111111101110110001011010010111000000111111011111111111111111111111111111111111111110110001101010011010111010111111001111010110110010,
	240'b101100011111111111100101110010101111111111111111111111111111111111111111111111111111111111110001101011101010011011100010111001111010101010101011111010011111111111111111111111111111111111111111111010011010101010111010111111001111010110110010,
	240'b101100011111111111100111101101101111011111111111111111111111111111111111111111111111111111110001101100001010100111100010111111011011110010100101110010011111111111111111111111111111111111111111111111001011110110111000111111001111010110110010,
	240'b101100011111111111101000101010111110001011111111111111111111111111111111111111111111111111110001101100001010100111100001111111111101101110100111101100001111000111111111111111111111111111111111111111111101100010111000111111001111010110110010,
	240'b101100011111111111101000101010011100010011111110111111111111111111111111111111111111111111110011101100001010100111100010111111111111100010110110101001101101001111111111111111111111111111111111111111111110111010111111111111001111010110110010,
	240'b101100001111111111101000101010101010110111101011111111111111111111111111111111111111100011100011101011111010100111010111111100001111000011000110101001101011011011111000111111111111111111111111111111111111101011001100111110101111010110110010,
	240'b101100001111111111101000101010111010011111000101111111101111111111111111111111111101010110101010101010101010101010101100101011101010111010101101101010011010111011110000111111111111111111111111111111111111111111011100111110101111010110110010,
	240'b101100001111111111101000101010111010100110101011111000101111111111111111111111111101000110100100101010101010101010100111101001101010011010100111101001101010101111101111111111111111111111111111111111111111111111101001111110111111010010110010,
	240'b101100001111111111101000101010111010101010101000101101111111010111111111111111111110010111000101101011001010101011000000110011011100110011001100110011001100111111110110111111111111111111111111111111111111111111110100111111001111010010110010,
	240'b101100001111111111101000101010111010101010101010101010001100011111111100111111111111111111110011101100001010100111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111011111010010110010,
	240'b101100001111111111101000101010111010101010101010101010101010100111010010111111101111111111110001101011111010100011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111011111010010110010,
	240'b101100011111111111101000101010111010101010101010101010101010100110101010110101001111111011111100111001011110001111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111011111010010110010,
	240'b101100011111111111101000101010111010101010101010101010101010101010101001101010101100111011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111001111010010110010,
	240'b101100011111111111101000101010111010101010101010101010101010101010101010101010011010100011000000111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111110101111010010110010,
	240'b101100011111111111101000101010111010101010101010101010101010100110101010101010101010101010101000101100001101000111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111000010111110111111010110110010,
	240'b101100011111111111101000101010111010100010100110101100011101100010110010101010011010101010101010101010011010100010110100110011101110101111111010111111111111111111111111111111111111111111111111111011111011101010111000111111001111010110110010,
	240'b101100001111111111101000101011101100000011000011110011111111101111001010101010101010101010101010101010101010101010101001101010001010110110111010110010111101100011100001111001011110010011010010101100111010011010111010111111001111010110110010,
	240'b101100001111111111100111101101001111001111111001111110001111111111101000101011011010100110101010101010101010101010101010101010101010100110101000101010001010100010101001101010111010101010101000101010011010100010111010111111001111010110110010,
	240'b101100001111111111100111101011101110101111011100110000101111011111000010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111001111010110110010,
	240'b101100001111111111101000101010011100110011101101101111011111011010111001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111001111010110110010,
	240'b101100001111111111101000101010101011000111110001110101001110000110110110101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111001111010110110010,
	240'b101100001111111111101000101010111010011111010111111010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111001111010110110010,
	240'b101010101111111111101011101011001010100010111000111101101100000010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111100111111101111000010101111,
	240'b100111011111111011111001101110101010011010101000110010101011111110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011111010010111111111101111110100001,
	240'b101101111110010111111111111011001100001010111001101110011011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100111011111001111111111100101110110011,
	240'b111100001011110011111000111111111111110111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111000111100011111110101,
	240'b111111101101100110111100111010101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011011010101111111111010011111110,
	240'b111100011111111011100110101010011010001010101010101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101011101010111010101110101011101010001001111010110010111010111111001111110010,
	240'b111110101111100011011110100101001001010110101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010001000110010110010111101011111101111111001,
	240'b111111111110100010111010110011001110000111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101101110011000101110100011111111111111110,
	240'b111110101011110011100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101101010111111110,
	240'b110010111101011111111111111011011001001001101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110101001101011011100111011001111111110111111011100010111001010,
	240'b101000001111101011111000010110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000010101000000000000100110100100111111111101100110100000,
	240'b101001011111111111001101000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101010101010000000010000000001000001111111011110110010101100,
	240'b101100001111111110111001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010011100011001011110000000000110000111101011111011010110010,
	240'b101100001111111110111001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000110100110111010100011010000000000110000111101011111011010110010,
	240'b101100001111111110111001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011001100110101010111110110010001010100101101111101011111011010110010,
	240'b101100001111111110111001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011101100111100010110110011100110101000101010111101011111011010110010,
	240'b101100001111111110111001000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110101101111010111000101111100111010110000110000111101001111011010110010,
	240'b101100011111111110111001000000110000000000001111010010010110011101100011010101000011001000010111000000000000000000000000000000000000000000000000000000000000000000010111101111101111000110011000100101000101110100110001111101001111011010110010,
	240'b101100011111111110111001000000000011101011000101111111001111111111111111111111101111011011010111101001010101110100011001000000000000000000000000000000000000000000000000010101111010110000000000000000000000000000110001111101011111011010110010,
	240'b101100011111111110110100001100001101111011111111111111111111111111111111111111111111111111111111111111111111111111011001011111010001100100000000000000000000000000000000000010000001000000000000000000000000000000110001111101011111011010110010,
	240'b101100011111111110111000101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001101010101000000010000000000000000000000000000000000000000000000000000000000110001111101011111011010110010,
	240'b101100011111111111010100111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100011100000110100000000000000000000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111111101010111101011111111111111111111111111111111111111111111111111111111111111111111110101110001011100000111101001111111111111111111111111010110000010101000000000000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111111101101111101101111111111111111111111111111111111111111111111111111111111111111111100110100110100011111011101101111111111111111111111111111111110110010000100110000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111111100111111100111111111111111111111111111111111111111111111111111111111111111111111111111000001100000000000101101101110011111111111111111111111111111111101000100000011100000000000000000000000000110001111101011111011010110010,
	240'b101100001111111111011101111011111111111111111111111111111111111111111111111111111111111111111111111111111101110100011001000000001000010111111111111111111111111111111111111111100111010100000000000000000000000000110001111101011111011010110010,
	240'b101100001111111111001100111001001111111111111111111111111111111111111111111111111111111111111111111111111111111101101010000000000010101111101101111111111111111111111111111111111110111000111000000000000000000000110001111101011111011010110010,
	240'b101100001111111111000000110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001000010100000000110100010111111111111111111111111111111111111111110110110000001110000000000110001111101011111011010110010,
	240'b101100011111111110110011100110001111111111111111111111111111111111111111111111111111111111101000011110100111000011001011010100010000000001000011111110001111111111111111111111111111111111111100010101000000000000110001111101011111011010110010,
	240'b101100011111111110110001011000001111111111111111111111111111111111111111111111111111111111010101000010110000000010101010101101100000001100000110101111011111111111111111111111111111111111111111101111000000010000101111111101011111011010110010,
	240'b101100011111111110110101001001001110011011111111111111111111111111111111111111111111111111010110000100100000000010100111111110000011010100000000010111011111111011111111111111111111111111111111111110000011100100101010111101011111011010110010,
	240'b101100011111111110111000000000111010100111111111111111111111111111111111111111111111111111010110000100100000000010100101111111111001001000000000000100101101010111111111111111111111111111111111111111111000100100101011111101011111011010110010,
	240'b101100011111111110111001000000000100110111111100111111111111111111111111111111111111111111011011000100100000000010101000111111111110100100100011000000000111101011111111111111111111111111111111111111111100110000111111111100101111011010110010,
	240'b101100001111111110111001000000010000101011000100111111111111111111111111111111111110100110101100000011110000000010000110110100111101001101010101000000000010010011101001111111111111111111111111111111111110111101100110111011111111011010110010,
	240'b101100001111111110111001000000110000000001010010111110111111111111111111111111111000000100001000000000010000000000000111000011000000110000001000000000000000101011010011111111111111111111111111111111111111110110010101111011011111011010110010,
	240'b101100001111111110111001000000110000000000000110101010011111111111111111111111110111010100000000000000000000000000000000000000000000000000000000000000000000001011010001111111111111111111111111111111111111111110111101111011111111011010110010,
	240'b101100001111111110111001000000110000000000000000001001111110000111111111111111111011000101010101000001110000000001000011011010010110011101100111011001100110110111100101111111111111111111111111111111111111111111011101111100111111010110110010,
	240'b101100001111111110111001000000110000000000000000000000000101011011110110111111111111111111011101000100100000000010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111101011111010110110010,
	240'b101100001111111110111001000000110000000000000000000000000000000001111000111111001111111111010110000011100000000010100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111101101111010110110010,
	240'b101100011111111110111001000000110000000000000000000000000000000000000010011111111111101111110101101100111010110111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101111111010110110010,
	240'b101100011111111110111001000000110000000000000000000000000000000000000000000000100110110011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110111101001111010110110010,
	240'b101100011111111110111001000000110000000000000000000000000000000000000000000000000000000001000010110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001111011101111011010110010,
	240'b101100011111111110111001000000110000000000000000000000000000000000000000000000000000000000000000000100110111010011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111100100101001000111100011111011010110010,
	240'b101100011111111110111001000000100000000000000000000101011000101000011001000000000000000000000000000000000000000000100000011011001100001011110001111111111111111111111111111111111111111111111111110100010011000100101011111101011111011010110010,
	240'b101100001111111110111000000010110100000101001101011011011111001101011111000000100000000000000000000000000000000000000000000000000000101000110001011000101000101110100110101100011010110101111000000111000000000000110001111101011111011010110010,
	240'b101100001111111110110110000111101101110011101110111010111111111110111010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111110111000000011001100010110010111010010011110100001001010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111110111001000000000110011011001010001110001110010000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111110111001000000010001010011010101011111011010010000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001111101011111011010110010,
	240'b101100001111111110111000000000110000000010000111110000000000110100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111101011111011010110010,
	240'b101010101111111111000001000001010000000000101001111001000100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101111110101111000110101111,
	240'b100111011111111011101100001011110000000000000000010111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111001111111111101111110100001,
	240'b101101111110010111111111110001100100101000101111001011000010111100110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100100110110111101101111111111100101110110011,
	240'b111100001011110011111000111111111111100111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011111111111111111111111000111100011111110101,
	240'b111111101101100110111100111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111011010101111111111010011111110,
	240'b111100011111111011100110101010011010001010101010101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101011101010111010101110101011101010001001111010110010111010111111001111110010,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule