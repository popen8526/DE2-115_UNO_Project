module green_six(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100001111011111110111101100111010001110101101101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011001001111110110101111100001111001011110010,
	240'b111011111111010011001111110001011101111011110000111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111011111101100110111110110011001111000011110001,
	240'b111011111100101011010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001011101001011101100,
	240'b110000001100010011111111111111011100011010100001101000001010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000001001111010011100101000101101000111111111111110101011111110111101,
	240'b100101001110000011111111101101110101010001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001001111010011110110100001110101010101010101101011001101111111111100101110100100,
	240'b101000111110110011111011011101110101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100110001111001011111010110010000101100110001100111111111101101110101111,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101101000011010001010000010111010111001011101111011111111111110011010111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010110111001001110011111110110011011011001111010111111111110011010111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101101101101111010111101100111111111011001101111010111111111110011010111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101101111100001000110101100001110111101011011101111010111111111110011010111011,
	240'b101100111111001111110101011010110101001001010100010100010100111101001111010100000101000101010010010101000101010101010101010101010101010101010101010101010101000101110100111100100111001101001101110011101011001001111010111111111110011010111011,
	240'b101100111111001111110101011010110100111101011011100001101010000010011111100101011000001001101010010110010101000001010010010101000101010101010101010101010101010001011100110101111101101010111100111101001000001001111100111111111110011010111011,
	240'b101100111111001111110101011010000110100111001100111110111111111111111111111111111111101011110000110100001010001101101111010101000101001001010101010101010101010101010010011101001100111011100010100111000101000101111111111111111110011010111011,
	240'b101100111111001111110011011101101101001011111111111111111111111111111111111111111111111111111111111111111111111111110000101111000111000101010001010101000101010101010101010100100101011001011001010100100100111110000000111111111110011010111011,
	240'b101100111111001111110000101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010011111010110000101001001010101010101010101010001010100010101010101000010000000111111111110011010111011,
	240'b101100111111001011110110111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000100110010001010001010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001011111101111101101111111111111111111111111111111111111111111111111111111111111111111111111111100111100111111010101111110111111111111111111101011001101001010100010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001011111110111110001111111111111111111111111111111111111111111111111111111111111111110001110111111001100101011010001000100011010110111111111111111111010111011001110101001001010101010101010101000010000000111111111110011010111011,
	240'b101100111111001011111100111100101111111111111111111111111111111111111111111111111111111010111000010110000100111001001110010011100100111001100001110011011111111111111111110010100101101101010011010101010101000010000000111111111110011010111011,
	240'b101100111111001011111000111001111111111111111111111111111111111111111111111111111110011001100010010011000101111110001011100001110101101001001111011100011111000011111111111111111010101101010010010101010101000010000000111111111110011010111011,
	240'b101100111111001111110010110110001111111111111111111111111111111111111111111111111111011110111000011101111100100011111110111111011011011101010110010100011100000011111111111111111111011101111111010100000101000010000000111111111110011010111011,
	240'b101100111111001111110000110000001111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111001111000010011001001111011111111111111111111111111010010010110100100111110000000111111111110011010111011,
	240'b101100111111001111110000100111101111110111111111111111111111111111111111111111111111111111111111111100111011101010010101100110001100001010000011010011001001001011111111111111111111111111111101100011110100101110000000111111111110011010111011,
	240'b101100111111001111110010100000001110110011111111111111111111111111111111111111111111111111100001011110100101000101001110010011100101010101011001010100001001001011111111111111111111111111111111110100100101001101111111111111111110011010111011,
	240'b101100111111001111110101011010111100011111111111111111111111111111111111111111111111001101111011010011100101001001100001010111100101000101010100010100001001001011111111111111111111111111111111111110100111100001111100111111111110011010111011,
	240'b101100111111001111110101011001101001001011111111111111111111111111111111111111111011110001010001010101001001101111100000110110111000101001010010010100001001001011111111111111111111111111111111111111111010101101111100111111111110011010111011,
	240'b101100111111001111110101011010010110000111100111111111111111111111111111111111101000111101001011011110101111100011111111111111111110101101101001010011011001001011111111111111111111111111111111111111111101011110000111111111111110011010111011,
	240'b101100111111001111110101011010110100111010100111111111111111111111111111111110110111111001001100100111111111111111111111111111111111111110000110010010111001001011111111111111111111111111111111111111111111000010011101111111111110011010111011,
	240'b101100111111001111110101011010110101000001100101111001101111111111111111111111011000010001001011100100001111111111111111111111111111101001111001010011001001110111111111111111111111111111111111111111111111110010111010111111011110011010111011,
	240'b101100111111001111110101011010110101001001010000100101011111110111111111111111111010010101001101011000001101000011111111111111101011110001010111010100001011111111111111111111111111111111111111111111111111111111010010111111101110011010111011,
	240'b101100111111001111110101011010110101001001010100010101111100010111111111111111111101111101100001010100000110001010010100100011010101110001001111011100001110111111111111111111111111111111111111111111111111111111100111111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010100100110100011011111111111111111111110110110010101100100111001001110010011100100111001011110110010111111111111111111111111111111111111111111111111111111111111110101111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010101010101000001111000111010011111111111111110110001000111111101101001011010101000011111010010111111111111111111111111111111111111111111111111111111111111111111111100111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010000011111011110011111111111111001001011000110100000101000011011011011101110111111111111111111111111111111111111111111111111111111111111111111111010111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010100000111001111011011110011001000011010001001100010001000011111011001111111111111111111111111111111111111111111111111111111111111111111100011111111101110010110111011,
	240'b101100111111001111110101011010110101001001010101010101000101010101010101010101010101000101100010101011101111010011111111111111101111110111111110111111111111111111111111111111111111111111111111111111111111100110110001111111101110011010111011,
	240'b101100111111001111110101011010110101000101010010010101110101001101010011010101010101010101010010010100110111110111000111111110001111111111111111111111111111111111111111111111111111111111111111111111111011110010000010111111111110011010111011,
	240'b101100111111001111110101011010100101011010100111110111111011110001100100010100110101010101010101010101010101000101010111011111001011010011011101111101111111111011111111111111111111111111111010110000110101111001111110111111111110011010111011,
	240'b101100111111001111110101011001111001100011110100101111011110100110111110010101000101010001010101010101010101010101010100010100010101000101011111011101001000110110100000101010011010010110000000010110000100111010000000111111111110011010111011,
	240'b101100111111001111110101011010101100110110110101010001111000111011101010011000110101001101010101010101010101010101010101010101010101010101010011010100010101000001001111010011110100111101010001010101000101000010000000111111111110011010111011,
	240'b101100111111001111110100011010111101010011000100010101101010001011100101010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001111110100011010111101000011111101111001011111010110100100010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001111110100011010111101000111001011101010101001000101010111010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001111110101011001111011011011011011011101001010101010001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001111111111111111110011010111011,
	240'b101000111110110011111010011100110110100111011101111110011110110110000111010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110001100111111111101101110110000,
	240'b100100101110000011111111101101000101000101011101011110100110011001001110010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011100101101011001010111111111100101110100011,
	240'b101111011100010111111111111111001100000010011010100110001001101010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111101100110011111111111110111011111110111010,
	240'b111011101100100011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001111101000011101010,
	240'b111110011111011011000101110001101110000111110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111100111101110111000100110100011111100111111001,
	240'b111111111111101111101001101010011001111010110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101011101001110110111110111111101111111111111110,
	240'b111100001111011111110111101100111010001110101101101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011001001111110110101111100001111001011110010,
	240'b111011111111010011001111110001011101111011110000111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111011111101100110111110110011001111000011110001,
	240'b111011111100101011010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001011101001011101100,
	240'b110000001100010011111110111111101110001011010000110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111011001110110100011110100011111111111110101011111110111101,
	240'b100101001110000011111111110110111010101010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111011010010111010101010101010110011100110111111111100101110100100,
	240'b101000111110110011111101101110111010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001110011001111100011111101111000111010110011000110111111111101101010101111,
	240'b101100111111001011111011101101011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110100001101000111000000111101011100101110111101111111111110011010111011,
	240'b101100111111001011111011101101011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011011100100111001111111011001101101010111101111111111110011010111011,
	240'b101100111111001011111011101101011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110110101111101011110101111111111101100110111100111111111110011010111011,
	240'b101100111111001011111011101101011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110110111110001100011010110000111011101101101110111100111111111110011010111011,
	240'b101100111111001011111011101101011010100110101001101010001010011110100111101001111010100010101001101010011010101010101010101010101010101010101010101010101010100010111001111110011011100110100110111001101101100110111101111111111110011010111011,
	240'b101100111111001011111011101101011010011110101101110000101101000011001111110010101100000010110101101011001010011110101000101010101010101010101010101010101010100110101110111010111110110011011101111110011100000010111101111111111110011010111011,
	240'b101100111111001011111011101100111011010011100110111111011111111111111111111111111111110111110111111010001101000110110111101010011010100010101010101010101010101010101001101110011110011011110001110011101010100010111111111111111110011010111011,
	240'b101100111111001011111010101110101110100111111111111111111111111111111111111111111111111111111111111111111111111111110111110111011011100010101000101010011010101010101010101010011010101110101100101010011010100010111111111111111110011010111011,
	240'b101100111111001011111000110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011001111101011001010100010101010101010101010101010101001101010101010100010111111111111111110011010111011,
	240'b101100111111001011111011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011001010101000101010101010101010101010101010101010100010111111111111111110011010111011,
	240'b101100111111000111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111110011110011111101011111111011111111111111111110101110110100101010001010101010101010101010101010100010111111111111111110011010111011,
	240'b101100111111000111111111111111001111111111111111111111111111111111111111111111111111111111111111111000111011111110110010101100111100001111101010111111111111111111101011101100111010100010101010101010101010100010111111111111111110011010111011,
	240'b101100111111000111111110111110001111111111111111111111111111111111111111111111111111111111011100101011001010011110100111101001101010011010110000111001101111111111111111111001011010110110101001101010101010100010111111111111111110011010111011,
	240'b101100111111001011111100111100111111111111111111111111111111111111111111111111111111001110110000101001101010111111000101110000111010110010100111101110001111011111111111111111111101010110101000101010101010100010111111111111111110011010111011,
	240'b101100111111001011111001111010111111111111111111111111111111111111111111111111111111101111011011101110111110001111111111111111101101101110101011101010001110000011111111111111111111101110111111101010001010100010111111111111111110011010111011,
	240'b101100111111001011111000111000001111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111010111100101001011100111011111111111111111111111111101000101011001010011110111111111111111110011010111011,
	240'b101100111111001011111001110011111111111011111111111111111111111111111111111111111111111111111111111110011101110011001010110011001110000111000001101001011100100011111111111111111111111111111110110001111010010110111111111111111110011010111011,
	240'b101100111111001011111010110000001111010111111111111111111111111111111111111111111111111111110000101111001010100010100110101001111010101010101100101001111100100011111111111111111111111111111111111010011010100110111111111111111110011010111011,
	240'b101100111111001011111011101101011110001111111111111111111111111111111111111111111111100110111101101001101010100110110000101011101010100010101010101001111100100011111111111111111111111111111111111111011011110010111101111111111110011010111011,
	240'b101100111111001011111011101100101100100011111111111111111111111111111111111111111101111010101000101010011100110111110000111011011100010010101001101001111100100011111111111111111111111111111111111111111101010110111101111111111110011010111011,
	240'b101100111111001011111011101101001011000011110011111111111111111111111111111111111100011110100101101111011111110011111111111111111111010110110100101001101100100011111111111111111111111111111111111111111110101111000011111111111110011010111011,
	240'b101100111111001011111011101101011010011011010011111111111111111111111111111111011011111110100101110011111111111111111111111111111111111111000011101001011100100011111111111111111111111111111111111111111111100011001110111111111110011010111011,
	240'b101100111111001011111011101101011010011110110010111100101111111111111111111111101100001010100101110001111111111111111111111111111111110110111100101001011100111011111111111111111111111111111111111111111111110111011100111111111110011010111011,
	240'b101100111111001011111011101101011010100110101000110010101111111011111111111111111101001010100110101011111110100011111111111111111101110110101011101010001101111111111111111111111111111111111111111111111111111111101001111111111110010110111011,
	240'b101100111111001011111011101101011010100110101001101010111110001011111111111111111110111110110000101001111011000111001010110001101010110110100111101101111111011111111111111111111111111111111111111111111111111111110011111111111110010110111011,
	240'b101100111111001011111011101101011010100110101010101010001011001111101111111111111111111111011011101010111010011110100111101001111010011110101111111001011111111111111111111111111111111111111111111111111111111111111001111111111110010110111011,
	240'b101100111111001011111011101101011010100110101010101010101010100010111011111101001111111111111111111000011011111110110100101101011100001111101000111111111111111111111111111111111111111111111111111111111111111111111101111111111110010110111011,
	240'b101100111111001011111011101101011010100110101010101010101010101010100111101111101111001111111111111100011101100011001111110100001101101011110110111111111111111111111111111111111111111111111111111111111111111111111101111111111110010110111011,
	240'b101100111111001011111011101101011010100110101010101010101010101010101010101010001011100111101101111001011100001111000100110001001100001111101100111111111111111111111111111111111111111111111111111111111111111111110001111111111110010110111011,
	240'b101100111111001011111011101101011010100110101010101010101010101010101010101010101010100010110001110101111111100111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111110011011000111111111110011010111011,
	240'b101100111111001011111011101101011010100010101001101010111010100110101001101010101010101010101001101010011011111011100011111111001111111111111111111111111111111111111111111111111111111111111111111111111101111011000000111111111110011010111011,
	240'b101100111111001011111011101101011010101111010011111011111101110110110010101010011010101010101010101010101010100010101011101111011101100111101110111110111111111111111111111111111111111111111101111000011010111010111110111111111110011010111011,
	240'b101100111111001011111011101100111100110011111001110111101111010011011111101010101010101010101010101010101010101010101010101010001010100010101111101110011100011011001111110101001101001011000000101010111010011110111111111111111110011010111011,
	240'b101100111111001011111011101101011110011011011010101000111100011111110100101100011010100110101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010101010100010111111111111111110011010111011,
	240'b101100111111001011111011101101011110100111100010101010111101000011110010101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111111111111111110011010111011,
	240'b101100111111001011111011101101011110011111111110111100101111101011010010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111111111111111110011010111011,
	240'b101100111111001011111011101101011110100011100110110101011100100010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111111111111111110011010111011,
	240'b101100111111001011111011101100111101101011101101101110101101010011000110101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111111111111111110011010111011,
	240'b101000111110110011111101101110011011010011101110111111001111011011000011101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111000101111111111101101110110000,
	240'b100100101110000011111111110110011010100010101110101111011011001110100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010110111100100111111111100101010100011,
	240'b101111011100010111111111111111101110000011001101110011001100110011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011111110011011111111111110111011111110111010,
	240'b111011101100100011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001111101000011101010,
	240'b111110011111011011000101110001101110000111110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111100111101110111000100110100011111100111111001,
	240'b111111111111101111101001101010011001111010110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101011101001110110111110111111101111111111111110,
	240'b111100001111011111110111101100111010001110101101101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011001001111110110101111100001111001011110010,
	240'b111011111111010011001111110001011101111011110000111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111011111101100110111110110011001111000011110001,
	240'b111011111100101011010010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001011101001011101100,
	240'b110000001100010011111111111111011100011010100001101000001010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000001001111010011100101000101101000111111111111110101011111110111101,
	240'b100101001110000011111111101101110101010001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001001111010011110110100001110101010101010101101011001101111111111100101110100100,
	240'b101000111110110011111011011101110101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100110001111001011111010110010000101100110001100111111111101101110101111,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101101000011010001010000010111010111001011101111011111111111110011010111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010110111001001110011111110110011011011001111010111111111110011010111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101101101101111010111101100111111111011001101111010111111111110011010111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101101111100001000110101100001110111101011011101111010111111111110011010111011,
	240'b101100111111001111110101011010110101001001010100010100010100111101001111010100000101000101010010010101000101010101010101010101010101010101010101010101010101000101110100111100100111001101001101110011101011001001111010111111111110011010111011,
	240'b101100111111001111110101011010110100111101011011100001101010000010011111100101011000001001101010010110010101000001010010010101000101010101010101010101010101010001011100110101111101101010111100111101001000001001111100111111111110011010111011,
	240'b101100111111001111110101011010000110100111001100111110111111111111111111111111111111101011110000110100001010001101101111010101000101001001010101010101010101010101010010011101001100111011100010100111000101000101111111111111111110011010111011,
	240'b101100111111001111110011011101101101001011111111111111111111111111111111111111111111111111111111111111111111111111110000101111000111000101010001010101000101010101010101010100100101011001011001010100100100111110000000111111111110011010111011,
	240'b101100111111001111110000101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010011111010110000101001001010101010101010101010001010100010101010101000010000000111111111110011010111011,
	240'b101100111111001011110110111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000100110010001010001010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001011111101111101101111111111111111111111111111111111111111111111111111111111111111111111111111100111100111111010101111110111111111111111111101011001101001010100010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001011111110111110001111111111111111111111111111111111111111111111111111111111111111110001110111111001100101011010001000100011010110111111111111111111010111011001110101001001010101010101010101000010000000111111111110011010111011,
	240'b101100111111001011111100111100101111111111111111111111111111111111111111111111111111111010111000010110000100111001001110010011100100111001100001110011011111111111111111110010100101101101010011010101010101000010000000111111111110011010111011,
	240'b101100111111001011111000111001111111111111111111111111111111111111111111111111111110011001100010010011000101111110001011100001110101101001001111011100011111000011111111111111111010101101010010010101010101000010000000111111111110011010111011,
	240'b101100111111001111110010110110001111111111111111111111111111111111111111111111111111011110111000011101111100100011111110111111011011011101010110010100011100000011111111111111111111011101111111010100000101000010000000111111111110011010111011,
	240'b101100111111001111110000110000001111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111001111000010011001001111011111111111111111111111111010010010110100100111110000000111111111110011010111011,
	240'b101100111111001111110000100111101111110111111111111111111111111111111111111111111111111111111111111100111011101010010101100110001100001010000011010011001001001011111111111111111111111111111101100011110100101110000000111111111110011010111011,
	240'b101100111111001111110010100000001110110011111111111111111111111111111111111111111111111111100001011110100101000101001110010011100101010101011001010100001001001011111111111111111111111111111111110100100101001101111111111111111110011010111011,
	240'b101100111111001111110101011010111100011111111111111111111111111111111111111111111111001101111011010011100101001001100001010111100101000101010100010100001001001011111111111111111111111111111111111110100111100001111100111111111110011010111011,
	240'b101100111111001111110101011001101001001011111111111111111111111111111111111111111011110001010001010101001001101111100000110110111000101001010010010100001001001011111111111111111111111111111111111111111010101101111100111111111110011010111011,
	240'b101100111111001111110101011010010110000111100111111111111111111111111111111111101000111101001011011110101111100011111111111111111110101101101001010011011001001011111111111111111111111111111111111111111101011110000111111111111110011010111011,
	240'b101100111111001111110101011010110100111010100111111111111111111111111111111110110111111001001100100111111111111111111111111111111111111110000110010010111001001011111111111111111111111111111111111111111111000010011101111111111110011010111011,
	240'b101100111111001111110101011010110101000001100101111001101111111111111111111111011000010001001011100100001111111111111111111111111111101001111001010011001001110111111111111111111111111111111111111111111111110010111010111111011110011010111011,
	240'b101100111111001111110101011010110101001001010000100101011111110111111111111111111010010101001101011000001101000011111111111111101011110001010111010100001011111111111111111111111111111111111111111111111111111111010010111111101110011010111011,
	240'b101100111111001111110101011010110101001001010100010101111100010111111111111111111101111101100001010100000110001010010100100011010101110001001111011100001110111111111111111111111111111111111111111111111111111111100111111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010100100110100011011111111111111111111110110110010101100100111001001110010011100100111001011110110010111111111111111111111111111111111111111111111111111111111111110101111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010101010101000001111000111010011111111111111110110001000111111101101001011010101000011111010010111111111111111111111111111111111111111111111111111111111111111111111100111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010000011111011110011111111111111001001011000110100000101000011011011011101110111111111111111111111111111111111111111111111111111111111111111111111010111111111110010110111011,
	240'b101100111111001111110101011010110101001001010101010101010101010101010101010100000111001111011011110011001000011010001001100010001000011111011001111111111111111111111111111111111111111111111111111111111111111111100011111111101110010110111011,
	240'b101100111111001111110101011010110101001001010101010101000101010101010101010101010101000101100010101011101111010011111111111111101111110111111110111111111111111111111111111111111111111111111111111111111111100110110001111111101110011010111011,
	240'b101100111111001111110101011010110101000101010010010101110101001101010011010101010101010101010010010100110111110111000111111110001111111111111111111111111111111111111111111111111111111111111111111111111011110010000010111111111110011010111011,
	240'b101100111111001111110101011010100101011010100111110111111011110001100100010100110101010101010101010101010101000101010111011111001011010011011101111101111111111011111111111111111111111111111010110000110101111001111110111111111110011010111011,
	240'b101100111111001111110101011001111001100011110100101111011110100110111110010101000101010001010101010101010101010101010100010100010101000101011111011101001000110110100000101010011010010110000000010110000100111010000000111111111110011010111011,
	240'b101100111111001111110101011010101100110110110101010001111000111011101010011000110101001101010101010101010101010101010101010101010101010101010011010100010101000001001111010011110100111101010001010101000101000010000000111111111110011010111011,
	240'b101100111111001111110100011010111101010011000100010101101010001011100101010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001111110100011010111101000011111101111001011111010110100100010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001111110100011010111101000111001011101010101001000101010111010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010000000111111111110011010111011,
	240'b101100111111001111110101011001111011011011011011011101001010101010001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001111111111111111110011010111011,
	240'b101000111110110011111010011100110110100111011101111110011110110110000111010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110001100111111111101101110110000,
	240'b100100101110000011111111101101000101000101011101011110100110011001001110010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011100101101011001010111111111100101110100011,
	240'b101111011100010111111111111111001100000010011010100110001001101010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111101100110011111111111110111011111110111010,
	240'b111011101100100011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001111101000011101010,
	240'b111110011111011011000101110001101110000111110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111100111101110111000100110100011111100111111001,
	240'b111111111111101111101001101010011001111010110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101011101001110110111110111111101111111111111110,
};
assign data = picture[addr];
endmodule