module green_nine(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100001111010111110100101011011001111010101001101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001110010100110111010001111001011110000,
	240'b111100001110101011000011110011111110101111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110101111001101101110111110100111110000,
	240'b111011101011110111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011110111101111,
	240'b101111011100111111111111111101011011000110010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101000111110001101100100001011001111110110111111111100110110111110,
	240'b100101111110111011111110100111100100111101001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001001111010011100110101110000100011001000100110110100001111111101111000110010001,
	240'b101010111111110011110000011001100101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100010011110111111111010111001100111010001100111111100011111100110100111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110111100000001110010110100111100010001100011111010011111101010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111010101000101001000010101000111101101001101001111010001111101010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100111111011011101001010001111111001001011100001100010111010011111101010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111010011110111011110100110011110110011101100001111010011111101010110111,
	240'b101110001111111111100111011000010101001101010011010100000100111101001111010100000101000101010010010100110101010101010101010101010101010101010101010101010101001101100011111001111010001001101000011101010101101001100100111010011111101010110111,
	240'b101110001111111111100111011000010100111101100001100100001010101110101000100111101000100101110001010111010101000101010001010101000101010101010101010101010101010101010100101110111110110010111100111010011000100101100000111010011111101010110111,
	240'b101110001111111111100111010111100111011011011010111111111111111111111111111111111111110111110101110110011010111001111000010101110101000101010100010101010101010101010011011000111011100011011110101010100101101101100011111010011111101010110111,
	240'b101110001111111111100100011101111110001111111111111111111111111111111111111111111111111111111111111111111111111111110110110010000111110101010011010100110101010101010101010100110101001101010111010100100101001001100100111010011111101010110111,
	240'b101110001111111111100100101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110001011000000101000101010101010101010101010101010100010101010101001101100100111010011111101010110111,
	240'b101110001111111111101111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000111000101010001010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111110110111111001111111111111111111111111111111111111111111111111111111111111111111111111111100011100101111001101111100111111111111111111110011101111011010100000101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111110110111110111111111111111111111111111111111111111111111111111111111111111111110001110111110101100100011001000111111011001001111111111111111111101000011110000101000001010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111110101111110101111111111111111111111111111111111111111111111111111111110110111010110000100111001001110010011100100111001011001101110101111111111111111111000010110101001010010010101010101001101100100111010011111101010110111,
	240'b101110001111111111110001111100001111111111111111111111111111111111111111111111111110000001100000010100000101111110001110100011010101111001001111011000101110001011111111111111111100100101011001010101000101001101100100111010011111101010110111,
	240'b101110001111111111101010110111101111111111111111111111111111111111111111111111111010011001001110010111011100100011111110111111101100010101011011010011101010100011111111111111111111111110011101010100000101001101100100111010011111101010110111,
	240'b101110001111111111100011110010001111111111111111111111111111111111111111111111101000001101001011100010101111111111111111111111111111111110000110010010111000011111111110111111111111111111101011011010110101000001100100111010011111101010110111,
	240'b101110001111111111100010101001011111111111111111111111111111111111111111111111000111100001001011100110111111111111111111111111111111111110010110010010111000000111111100111111111111111111111111101100100100111101100100111010011111101010110111,
	240'b101110001111111111100011100000101111010111111111111111111111111111111111111111000111100001001101011110011111011111111111111111111111011001110110010011001001000011111111111111111111111111111111111011010110100001100001111010011111101010110111,
	240'b101110001111111111100110011001101101011011111111111111111111111111111111111111000111100001010001010101001001101111100101111001001001100101010011010100011011111011111111111111111111111111111111111111111001111001011111111010011111101010110111,
	240'b101110001111111111100111010111001010001011111111111111111111111111111111111111000111100001010001010101000101001001100100011000110101001001001110011111001111001111111111111111111111111111111111111111111101001001100111111010001111101010110111,
	240'b101110001111111111100111010111100110101011110000111111111111111111111111111111000111100001010001010110000101001001001110010011100101000001110111111000011111111111111111111111111111111111111111111111111111001110000001111001101111101010110111,
	240'b101110001111111111100111011000010101000010110101111111111111111111111111111111000111100001001101100100001011011010001110100100101011011011110001111111111111111111111111111111111111111111111111111111111111111110100011111001001111101010110111,
	240'b101110001111111111100111011000010100111101101101111011101111111111111111111111101000001101001011100011011111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111000101111001101111101010110111,
	240'b101110001111111111100111011000010101001101010001101000001111111111111111111111111010010001001101010111101100110111111111111111111100010110000000110001101111101011111111111111111111111111111111111111111111111111011111111010011111100110110111,
	240'b101110001111111111100111011000010101001101010011010110111100111011111111111111111101111001100000010100000110001010010101100100110101111101001100011001011110100111111111111111111111111111111111111111111111111111101011111100001111100010110111,
	240'b101110001111111111100111011000010101001101010101010100010110111011100101111111111111111110110100010101100100111001001110010011110100111101010111101101011111111011111111111111111111111111111111111111111111111111110001111101011111100010110111,
	240'b101110001111111111100111011000010101001101010101010101010101000001111110111011011111111111111110110000100111110101100110011001010111110111000100111111101111111111111111111111111111111111111111111111111111111111110101111110001111100010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010000100000101110101011111111111010001011011010100010101000011011011011101010111111111111111111111111111111111111111111111111111111111111111111110100111101111111100010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010100000111011111011110110011011000000110000101100001011000000011001100111111111111111111111111111111111111111111111111111111111111111111101010111011111111100010110111,
	240'b101110001111111111100111011000010101001101010101010101000101010101010101010101010101000101100101101100101111001111111110111111001111101011111101111111111111111111111111111111111111111111111111111111111111111110111110111001101111101010110111,
	240'b101110001111111111100111011000010101001001010001010101000101001001010011010101010101010101010010010101001000000011001001111110101111111111111111111111111111111111111111111111111111111111111111111111111110000101111000111001111111101010110111,
	240'b101110001111111111100111011000000101101110100110110101111011000001011111010100110101010101010101010101000101000001011000011111101011011111100000111110011111111111111111111111111111111111111111110111010111100001100000111010011111101010110111,
	240'b101110001111111111100111010111011000110111101101110001001110111110110011010100110101010101010101010101010101010101010100010100010101001001100000011110001001001010100111101100011011001010010011011000100100111101100100111010011111101010110111,
	240'b101110001111111111100111011000010101110001110110011000111010001111101000010111100101001101010101010101010101010101010101010101010101010101010011010100010101000001010000010100000101000001010000010100110101001101100100111010011111101010110111,
	240'b101110001111111111100111010111110110011011001100111100101110101011101100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111100110010111111011101011100100100101101101100011101110011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111100110011001011110000010011110010000101000110111101110011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111100110011000001100101111001100011010111011111011011010010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101010111111110011101111011000100111101111101011111101111111000010001010010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101010111100001111100110101000,
	240'b100101101110111111111110100110100100110001101001100010000110111101001110010011110101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110100111110011110111111101111000110010000,
	240'b101110011101000111111111111101001010101110001010100010011000101110001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011011010110111110101111111111100111110111010,
	240'b111011011011101111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101011101111101101,
	240'b111110001110111010111101110100101110111011111100111111011111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111101111111001110110111010010110000001110111111111000,
	240'b111111111111111111100110101000111001101010110000101100111011001110110011101100111011001110110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110011101011111001101010101101111101101111111111111111,
	240'b111100001111010111110100101011011001111010101001101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001110010100110111010001111001011110000,
	240'b111100001110101011000011110011111110101111111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001110101111001101101110111110100111110000,
	240'b111011101011110111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011110111101111,
	240'b101111011100111111111111111110101101100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100011111000110110001111101100111111011111111111100110110111110,
	240'b100101111110111011111111110011111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001101011010111000001101100011010011011010000111111111111000010010001,
	240'b101010111111101111111000101100111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110001001111011111111101111100111011101010110011111110001111011110100111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101101111011011101111110111000111010011110001010110001111101001111100010110111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110011111101011100010010100001110100011110110010110100111101001111100010110111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110011111101101110100011000111111100011101110010110000111101011111100010110111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110011111101001111011111111010111001111011001110110000111101011111100010110111,
	240'b101110001111111111110011101100001010100110101001101010001010011110100111101001111010100010101000101010011010101010101010101010101010101010101010101010101010100110110001111100111101000110110011101110101010110010110001111101011111100010110111,
	240'b101110001111111111110011101100001010011110110000110010001101010111010100110011101100010010111000101011101010100010101000101010101010101010101010101010101010101010101001110111011111010111011101111101001100010010101111111101011111100010110111,
	240'b101110001111111111110011101011101011101111101100111111111111111111111111111111111111111011111010111011001101011110111100101010111010100010101010101010101010101010101001101100011101101111101111110101001010110110110001111101011111100010110111,
	240'b101110001111111111110001101110111111000111111111111111111111111111111111111111111111111111111111111111111111111111111010111001001011111010101001101010011010101010101010101010011010100110101011101010011010100010110010111101011111100010110111,
	240'b101110001111111111110001110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011011000101011111010100010101010101010101010101010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111110111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011011100010101000101010101010101010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111111010111111011111111111111111111111111111111111111111111111111111111111111111111111111111110011110010111100101111110011111111111111111111001110111101101010001010101010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111111010111111011111111111111111111111111111111111111111111111111111111111111111111000111011111010110001101100011011111011100100111111111111111111110100101111001010100010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111111010111111011111111111111111111111111111111111111111111111111111111111011011101011001010011110100111101001111010011110101100110111011111111111111111111100001011010110101000101010101010100110110010111101011111100010110111,
	240'b101110001111111111111000111101111111111111111111111111111111111111111111111111111110111110110000101001111010111111000111110001101010111110100111101100011111000011111111111111111110010010101100101010011010100110110010111101011111100010110111,
	240'b101110001111111111110101111011101111111111111111111111111111111111111111111111111101001010100110101011101110010011111111111111111110001010101101101001111101010011111111111111111111111111001110101010001010100110110010111101011111100010110111,
	240'b101110001111111111110001111000111111111111111111111111111111111111111111111111101100000110100101110001001111111111111111111111111111111111000011101001011100001111111110111111111111111111110101101101011010011110110010111101011111100010110111,
	240'b101110001111111111110000110100101111111111111111111111111111111111111111111111011011110010100101110011011111111111111111111111111111111111001010101001011100000011111101111111111111111111111111110110001010011110110010111101011111100010110111,
	240'b101110001111111111110001110000011111101011111111111111111111111111111111111111011011101110100110101111001111101111111111111111111111101010111010101001011100100011111111111111111111111111111111111101101011001110110000111101011111100010110111,
	240'b101110001111111111110010101100101110101011111111111111111111111111111111111111011011101110101000101010101100110111110010111100101100110010101001101010001101111011111111111111111111111111111111111111111100111010101111111101011111100010110111,
	240'b101110001111111111110011101011101101000111111111111111111111111111111111111111011011101110101000101010011010100110110001101100011010100110100110101111011111100111111111111111111111111111111111111111111110100010110011111101001111100010110111,
	240'b101110001111111111110011101011111011010111110111111111111111111111111111111111011011101110101000101011001010100110100110101001101010100010111011111100001111111111111111111111111111111111111111111111111111100111000000111100111111100010110111,
	240'b101110001111111111110011101100001010100011011010111111111111111111111111111111011011101110100110110001111101101011000110110010001101101011111000111111111111111111111111111111111111111111111111111111111111111111010001111100101111100010110111,
	240'b101110001111111111110011101100001010011110110110111101101111111111111111111111101100000110100101110001101111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111100010111100111111100010110111,
	240'b101110001111111111110011101100001010100110101000110011111111111111111111111111111101000110100110101011111110011011111111111111111110001011000000111000101111110011111111111111111111111111111111111111111111111111101111111101001111100010110111,
	240'b101110001111111111110011101100001010100110101001101011011110011111111111111111111110111010101111101001111011000011001010110010011010111110100110101100101111010011111111111111111111111111111111111111111111111111110101111110001111100010110111,
	240'b101110001111111111110011101100001010100110101010101010001011011011110010111111111111111111011010101010111010011110100111101001111010011110101011110110101111111111111111111111111111111111111111111111111111111111111000111110101111011110110111,
	240'b101110001111111111110011101100001010100110101010101010101010100010111111111101101111111111111110111000001011111010110011101100101011111011100001111111111111111111111111111111111111111111111111111111111111111111111010111111001111011110110111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101000110000001111010111111111111101001101101011010000110100001101101011110100111111111111111111111111111111111111111111111111111111111111111111111010111111001111011110110111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101010101010001011101111101111111001101100000011000010110000101011111111100110111111111111111111111111111111111111111111111111111111111111111111110101111101111111100010110111,
	240'b101110001111111111110011101100001010100110101010101010101010101010101010101010101010100010110010110110011111100111111111111111011111110111111110111111111111111111111111111111111111111111111111111111111111111111011111111100111111100010110111,
	240'b101110001111111111110011101100001010100010101000101010101010100010101001101010101010101010101001101010101011111111100100111111001111111111111111111111111111111111111111111111111111111111111111111111111111000010111100111100111111100010110111,
	240'b101110001111111111110011101100001010110111010010111010111101011110101111101010011010101010101010101010101010100010101011101111111101101111101111111111001111111111111111111111111111111111111111111011101011101110110000111101011111100010110111,
	240'b101110001111111111110011101011101100011011110110111000011111011111011001101010011010101010101010101010101010101010101001101010001010100010110000101110111100100011010011110110001101100011001001101100001010011110110010111101011111100010110111,
	240'b101110001111111111110011101100001010111010111010101100011101000111110011101011101010100110101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100110110010111101011111100010110111,
	240'b101110001111111111110011101011111011001111100101111110001111010011110101101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111110011101011111101110111110010110010111110110011110111101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111110010101100101111000011001111101000001100011011110111101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101011111100010110111,
	240'b101110001111111111110011101100001110010111100101101101011101111111101101101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101011111100010110111,
	240'b101010111111101111111000101100011011110111110101111110111111100011000100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110100111110001111011110101000,
	240'b100101101110111111111111110011011010011010110100110001001011011110100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011111001110111111111111000110010000,
	240'b101110011101000111111111111110011101010111000101110001001100010111000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101101011011111010111111111100111110111010,
	240'b111011011011101111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101011101111101101,
	240'b111110001110111010111101110100101110111011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001110110111010010110000001110111111111000,
	240'b111111111111111111100110101000111001101010110000101100111011001110110011101100111011001110110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110011101011111001101010101101111101101111111111111111,
	240'b111100001111010111110100101011011001111010101001101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101010101010111010101110101011101010011001110010100110111010001111001011110000,
	240'b111100001110101011000011110011111110101111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110101111001101101110111110100111110000,
	240'b111011101011110111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011110111101111,
	240'b101111011100111111111111111101011011000110010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101000111110001101100100001011001111110110111111111100110110111110,
	240'b100101111110111011111110100111100100111101001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001001111010011100110101110000100011001000100110110100001111111101111000110010001,
	240'b101010111111110011110000011001100101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100010011110111111111010111001100111010001100111111100011111100110100111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110111100000001110010110100111100010001100011111010011111101010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111010101000101001000010101000111101101001101001111010001111101010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100111111011011101001010001111111001001011100001100010111010011111101010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101000111010011110111011110100110011110110011101100001111010011111101010110111,
	240'b101110001111111111100111011000010101001101010011010100000100111101001111010100000101000101010010010100110101010101010101010101010101010101010101010101010101001101100011111001111010001001101000011101010101101001100100111010011111101010110111,
	240'b101110001111111111100111011000010100111101100001100100001010101110101000100111101000100101110001010111010101000101010001010101000101010101010101010101010101010101010100101110111110110010111100111010011000100101100000111010011111101010110111,
	240'b101110001111111111100111010111100111011011011010111111111111111111111111111111111111110111110101110110011010111001111000010101110101000101010100010101010101010101010011011000111011100011011110101010100101101101100011111010011111101010110111,
	240'b101110001111111111100100011101111110001111111111111111111111111111111111111111111111111111111111111111111111111111110110110010000111110101010011010100110101010101010101010100110101001101010111010100100101001001100100111010011111101010110111,
	240'b101110001111111111100100101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110001011000000101000101010101010101010101010101010100010101010101001101100100111010011111101010110111,
	240'b101110001111111111101111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000111000101010001010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111110110111111001111111111111111111111111111111111111111111111111111111111111111111111111111100011100101111001101111100111111111111111111110011101111011010100000101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111110110111110111111111111111111111111111111111111111111111111111111111111111111110001110111110101100100011001000111111011001001111111111111111111101000011110000101000001010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111110101111110101111111111111111111111111111111111111111111111111111111110110111010110000100111001001110010011100100111001011001101110101111111111111111111000010110101001010010010101010101001101100100111010011111101010110111,
	240'b101110001111111111110001111100001111111111111111111111111111111111111111111111111110000001100000010100000101111110001110100011010101111001001111011000101110001011111111111111111100100101011001010101000101001101100100111010011111101010110111,
	240'b101110001111111111101010110111101111111111111111111111111111111111111111111111111010011001001110010111011100100011111110111111101100010101011011010011101010100011111111111111111111111110011101010100000101001101100100111010011111101010110111,
	240'b101110001111111111100011110010001111111111111111111111111111111111111111111111101000001101001011100010101111111111111111111111111111111110000110010010111000011111111110111111111111111111101011011010110101000001100100111010011111101010110111,
	240'b101110001111111111100010101001011111111111111111111111111111111111111111111111000111100001001011100110111111111111111111111111111111111110010110010010111000000111111100111111111111111111111111101100100100111101100100111010011111101010110111,
	240'b101110001111111111100011100000101111010111111111111111111111111111111111111111000111100001001101011110011111011111111111111111111111011001110110010011001001000011111111111111111111111111111111111011010110100001100001111010011111101010110111,
	240'b101110001111111111100110011001101101011011111111111111111111111111111111111111000111100001010001010101001001101111100101111001001001100101010011010100011011111011111111111111111111111111111111111111111001111001011111111010011111101010110111,
	240'b101110001111111111100111010111001010001011111111111111111111111111111111111111000111100001010001010101000101001001100100011000110101001001001110011111001111001111111111111111111111111111111111111111111101001001100111111010001111101010110111,
	240'b101110001111111111100111010111100110101011110000111111111111111111111111111111000111100001010001010110000101001001001110010011100101000001110111111000011111111111111111111111111111111111111111111111111111001110000001111001101111101010110111,
	240'b101110001111111111100111011000010101000010110101111111111111111111111111111111000111100001001101100100001011011010001110100100101011011011110001111111111111111111111111111111111111111111111111111111111111111110100011111001001111101010110111,
	240'b101110001111111111100111011000010100111101101101111011101111111111111111111111101000001101001011100011011111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111000101111001101111101010110111,
	240'b101110001111111111100111011000010101001101010001101000001111111111111111111111111010010001001101010111101100110111111111111111111100010110000000110001101111101011111111111111111111111111111111111111111111111111011111111010011111100110110111,
	240'b101110001111111111100111011000010101001101010011010110111100111011111111111111111101111001100000010100000110001010010101100100110101111101001100011001011110100111111111111111111111111111111111111111111111111111101011111100001111100010110111,
	240'b101110001111111111100111011000010101001101010101010100010110111011100101111111111111111110110100010101100100111001001110010011110100111101010111101101011111111011111111111111111111111111111111111111111111111111110001111101011111100010110111,
	240'b101110001111111111100111011000010101001101010101010101010101000001111110111011011111111111111110110000100111110101100110011001010111110111000100111111101111111111111111111111111111111111111111111111111111111111110101111110001111100010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010000100000101110101011111111111010001011011010100010101000011011011011101010111111111111111111111111111111111111111111111111111111111111111111110100111101111111100010110111,
	240'b101110001111111111100111011000010101001101010101010101010101010101010101010100000111011111011110110011011000000110000101100001011000000011001100111111111111111111111111111111111111111111111111111111111111111111101010111011111111100010110111,
	240'b101110001111111111100111011000010101001101010101010101000101010101010101010101010101000101100101101100101111001111111110111111001111101011111101111111111111111111111111111111111111111111111111111111111111111110111110111001101111101010110111,
	240'b101110001111111111100111011000010101001001010001010101000101001001010011010101010101010101010010010101001000000011001001111110101111111111111111111111111111111111111111111111111111111111111111111111111110000101111000111001111111101010110111,
	240'b101110001111111111100111011000000101101110100110110101111011000001011111010100110101010101010101010101000101000001011000011111101011011111100000111110011111111111111111111111111111111111111111110111010111100001100000111010011111101010110111,
	240'b101110001111111111100111010111011000110111101101110001001110111110110011010100110101010101010101010101010101010101010100010100010101001001100000011110001001001010100111101100011011001010010011011000100100111101100100111010011111101010110111,
	240'b101110001111111111100111011000010101110001110110011000111010001111101000010111100101001101010101010101010101010101010101010101010101010101010011010100010101000001010000010100000101000001010000010100110101001101100100111010011111101010110111,
	240'b101110001111111111100111010111110110011011001100111100101110101011101100011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111100110010111111011101011100100100101101101100011101110011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111100110011001011110000010011110010000101000110111101110011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101110001111111111100110011000001100101111001100011010111011111011011010010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010011111101010110111,
	240'b101010111111110011101111011000100111101111101011111101111111000010001010010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101010111100001111100110101000,
	240'b100101101110111111111110100110100100110001101001100010000110111101001110010011110101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110100111110011110111111101111000110010000,
	240'b101110011101000111111111111101001010101110001010100010011000101110001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011011010110111110101111111111100111110111010,
	240'b111011011011101111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101011101111101101,
	240'b111110001110111010111101110100101110111011111100111111011111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111101111111001110110111010010110000001110111111111000,
	240'b111111111111111111100110101000111001101010110000101100111011001110110011101100111011001110110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110011101011111001101010101101111101101111111111111111,
};
assign data = picture[addr];
endmodule