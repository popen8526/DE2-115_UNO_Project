module red_seven(
    input [7:0] addr,
    output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111011111111011111101000101111101011000010110010101100101011001010110010101100101011001010110011101100111011001110110011101100111011001010110010101100101011001010110010101100111011001110110011101100101011000010111110111001001111000111101111,
	240'b111100101101111110111111111000101111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100011011100101110001101111011110010,
	240'b111000101011110011110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011101011101000,
	240'b101101001110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110110101,
	240'b100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010001111,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110100101,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b101110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110101101,
	240'b101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010010100,
	240'b101001001111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010011111,
	240'b110100011100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000111011000,
	240'b111100001100100011010001111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110001111100100111110001,
	240'b111101101111011111001001101011101011101011000100110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100010110000110100001111011111110110,
	240'b111011111111011111101000101111101011000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011000110111111111001001111001011101111,
	240'b111100101101111110111111111000101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111100011011100101110001101111011110010,
	240'b111000101011110011110101111111111111111111111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110111111111111111111111011111011101011101000,
	240'b101101001110010111111111111000101001011101111110011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011110110111101001111010011110111001100111101010111111111101101110110101,
	240'b100110111111111111110100011110110100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001011000100100011001111010011110100111011000110010001111111110101111101110001111,
	240'b101100101111111111010100010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010101111000111100111111100101110100001101001111000101111111110100101,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101011011010001011110100110011110100001100101110111001111111110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000101000001101100101010110011001111000101001011110110111011111111110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011011101110101001111101010011110101000001011010110111101111111110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101011100110010110011010100000101010001011010110111101111111110110001,
	240'b101111001111111111001101010100110101010101010011010100000101000101010001010100000101000001010010010101000101010101010101010101010101010101010101010101010101010101010101010100001001010111100001010111110101001001011010110111101111111110110001,
	240'b101111001111111111001101010100100101000101101000100101101010100110100111100111101000101101110011010110110101000101010001010101000101010101010101010101010101010101010101010100110110011111101010100010100100111101011010110111101111111110110001,
	240'b101111001111111111001101010011111000101011100100111111111111111111111111111111111111111011110010110110011010110101111000010101010101000101010101010101010101010101010101010101010101010010101111100111110101000101011001110111101111111110110001,
	240'b101111001111111111001001011110111111001011111111111111111111111111111111111111111111111111111111111111111111111111110100110000010111100001010010010100110101010101010101010101010101010101011000010110100101010001011010110111101111111110110001,
	240'b101111001111111111001111110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101010010111100101000101010101010101010101010101010100010101000101010001011010110111101111111110110001,
	240'b101111001111111111101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000110111101010000010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111111011111111001111111111111111111111111111111111111111111011111110010111100110111001101110011011100110111001101110011011100110111011001101111101111001010100000101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111111100111111011111111111111111111111111111111111111111100110000101111001100010011000100110001001100010011000100110001001100000011011001110101111101000011101010101000101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111111000111110101111111111111111111111111111111111111111100011010100111001010010010011100100111001001110010011100101000001010001010111011110010011111111110111100110011101010010010101010101010001011010110111101111111110110001,
	240'b101111001111111111101111111101001111111111111111111111111111111111111111100100100100111101100000100010011000101010001010100010110111011101010010010111111110010011111111111111111100010001011000010101000101010001011010110111101111111110110001,
	240'b101111001111111111100000111010101111111111111111111111111111111111111111101110010101000001100101111010011111111111111111111111111100001001010001010111111110010011111111111111111111111010011010010100000101010001011010110111101111111110110001,
	240'b101111001111111111010011110110101111111111111111111111111111111111111111111010000110010001010000101110101111111111111111111111111011111101001011010110101110001111111111111111111111111111101010011010100101000101011010110111101111111110110001,
	240'b101111001111111111001011101110101111111111111111111111111111111111111111111111101000111101001011100001001111110011111111111111111110010010110011101110011111001111111111111111111111111111111111101100100101000101011001110111101111111110110001,
	240'b101111001111111111001000100101101111111111111111111111111111111111111111111111111100010001010010010111101110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111011100110101001010111110111101111111110110001,
	240'b101111001111111111001010011011001111001011111111111111111111111111111111111111111110111001101010010011101010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001001010101110111101111111110110001,
	240'b101111001111111111001100010101001100101111111111111111111111111111111111111111111111111110011000010010110111101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111101011101011111110111011111111110110001,
	240'b101111001111111111001101010011101000111011111110111111111111111111111111111111111111111111001101010101010101101011011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111101110110101111111110110001,
	240'b101111001111111111001101010100010101111011011101111111111111111111111111111111111111111111110100011100010100110010100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001110110001111111110110001,
	240'b101111001111111111001101010100100101000010010010111111101111111111111111111111111111111111111111101000100100110001110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111000101110110111111111010110001,
	240'b101111001111111111001101010100110101001101011010110011011111111111111111111111111111111111111111110101100101100001010101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111000011111111010110001,
	240'b101111001111111111001101010100110101010101010001011101001111000011111111111111111111111111111111111110000111100101001100100110101111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111011011111110110110001,
	240'b101111001111111111001101010100110101010101010101010100011001010111111011111111111111111111111111111111111010110001001101011010111111000011111111111111111111111111111111111111111111111111111111111111111111111111110100111101011111110010110001,
	240'b101111001111111111001101010100110101010101010101010101000101001110101011111111101111111111111111111111111101111101011011010011111100001111111111111111111111111111111111111111111111111111111111111111111111111111111000111110011111101110110001,
	240'b101111001111111111001101010100110101010101010101010101010101001101010111101100001111111011111111111111111111101111000001101100001101011011111111111111111111111111111111111111111111111111111111111111111111111111111010111110111111101110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010011010101111010010111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111110010110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010100110101001110001101111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111000011111111010110001,
	240'b101111001111111111001101010100110101010101010010010100100101010101010101010101010101010001010000011010101011010111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010010110110011111111110110001,
	240'b101111001111111111001101010100100101010110001110011111000101001001010101010101010101010101010101010100100101001101110110101100111110011011111110111111111111111111111111111111111111111111111111111110111010101001011010110111011111111110110001,
	240'b101111001111111111001101010100100101000010110010110100010101010101010100010101010101010101010101010101010101010101010001010100100110011010000111101011101100100111011001111000011110001011001100100011010101010001011001110111101111111110110001,
	240'b101111001111111111001101010100110101000101111001111011000111001001010010010101010101010101010101010101010101010101010101010101010101001101010001010100000101010001011101011000110110001101010111010100010101001101011010110111101111111110110001,
	240'b101111001111111111001101010100110101001101011000110110001010010101010000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010011010100110101001101010100010101010101010001011010110111101111111110110001,
	240'b101111001111111111001101010100110101001001001111101001001101100001011001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111001101010101010110001001010100011100001110101101111010010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111001010011001101101100001110001010100001100110110110000010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101110001111111111001100011010101111100111001011101101101110000111011011010110000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111111111111110101101,
	240'b101000011111111111100100011101001100100011011001110110101101100110111000010110000101001101010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000100111101101111111100011111111010010100,
	240'b101001001111010011111111101110010110100001011101010111100101111001011101010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110010110100111000111111111111110110010011111,
	240'b110100011100100111111111111111111110010111010111110110001101100011011000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011110100111111111111111101100000111011000,
	240'b111100001100100011010001111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110001111100100111110001,
	240'b111101101111011111001001101011101011101011000100110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100010110000110100001111011111110110,
	240'b111011111111011111101000101111101011000010110010101100101011001010110010101100101011001010110011101100111011001110110011101100111011001010110010101100101011001010110010101100111011001110110011101100101011000010111110111001001111000111101111,
	240'b111100101101111110111111111000101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111100111011100101110001101111011110010,
	240'b111000101011110011110101111111111111111111111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110111111111111111111111011111011101011101000,
	240'b101101001110010111111111111000101001011101111110011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011110110111101001111010011110111001100111101010111111111101101110110101,
	240'b100110111111111111110100011110110100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001011000100100011001111010011110100111011000110010001111111110101111101110001111,
	240'b101100101111111111010100010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100100111010101111000111100111111100101110100001101001111000101111111110100101,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110101011011010001011110100110011110100001100101110111001111111110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000101000001101100101010110011001111000101001011110110111011111111110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011011101110101001111101010011110101000001011010110111101111111110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101011100110010110011010100000101010001011010110111101111111110110001,
	240'b101111001111111111001101010100110101010101010011010100000101000101010001010100000101000001010010010101000101010101010101010101010101010101010101010101010101010101010101010100001001010111100001010111110101001001011010110111101111111110110001,
	240'b101111001111111111001101010100100101000101101000100101101010100110100111100111101000101101110011010110110101000101010001010101000101010101010101010101010101010101010101010100110110011111101010100010100100111101011010110111101111111110110001,
	240'b101111001111111111001101010011111000101011100100111111111111111111111111111111111111111011110010110110011010110101111000010101010101000101010101010101010101010101010101010101010101010010101111100111110101000101011001110111101111111110110001,
	240'b101111001111111111001001011110111111001011111111111111111111111111111111111111111111111111111111111111111111111111110100110000010111100001010010010100110101010101010101010101010101010101011000010110100101010001011010110111101111111110110001,
	240'b101111001111111111001111110010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101010010111100101000101010101010101010101010101010100010101000101010001011010110111101111111110110001,
	240'b101111001111111111101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000110111101010000010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111111011111111001111111111111111111111111111111111111111111011111110010111100110111001101110011011100110111001101110011011100110111011001101111101111001010100000101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111111100111111011111111111111111111111111111111111111111100110000101111001100010011000100110001001100010011000100110001001100000011011001110101111101000011101010101000101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111111000111110101111111111111111111111111111111111111111100011010100111001010010010011100100111001001110010011100101000001010001010111011110010011111111110111100110011101010010010101010101010001011010110111101111111110110001,
	240'b101111001111111111101111111101001111111111111111111111111111111111111111100100100100111101100000100010011000101010001010100010110111011101010010010111111110010011111111111111111100010001011000010101000101010001011010110111101111111110110001,
	240'b101111001111111111100000111010101111111111111111111111111111111111111111101110010101000001100101111010011111111111111111111111111100001001010001010111111110010011111111111111111111111010011010010100000101010001011010110111101111111110110001,
	240'b101111001111111111010011110110101111111111111111111111111111111111111111111010000110010001010000101110101111111111111111111111111011111101001011010110101110001111111111111111111111111111101010011010100101000101011010110111101111111110110001,
	240'b101111001111111111001011101110101111111111111111111111111111111111111111111111101000111101001011100001001111110011111111111111111110010010110011101110011111001111111111111111111111111111111111101100100101000101011001110111101111111110110001,
	240'b101111001111111111001000100101101111111111111111111111111111111111111111111111111100010001010010010111101110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111011100110101001010111110111101111111110110001,
	240'b101111001111111111001010011011001111001011111111111111111111111111111111111111111110111001101010010011101010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001001010101110111101111111110110001,
	240'b101111001111111111001100010101001100101111111111111111111111111111111111111111111111111110011000010010110111101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111101011101011111110111011111111110110001,
	240'b101111001111111111001101010011101000111011111110111111111111111111111111111111111111111111001101010101010101101011011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111101110110101111111110110001,
	240'b101111001111111111001101010100010101111011011101111111111111111111111111111111111111111111110100011100010100110010100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001110110001111111110110001,
	240'b101111001111111111001101010100100101000010010010111111101111111111111111111111111111111111111111101000100100110001110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111000101110110111111111010110001,
	240'b101111001111111111001101010100110101001101011010110011011111111111111111111111111111111111111111110101100101100001010101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111000011111111010110001,
	240'b101111001111111111001101010100110101010101010001011101001111000011111111111111111111111111111111111110000111100101001100100110101111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111011011111110110110001,
	240'b101111001111111111001101010100110101010101010101010100011001010111111011111111111111111111111111111111111010110001001101011010111111000011111111111111111111111111111111111111111111111111111111111111111111111111110100111101011111110010110001,
	240'b101111001111111111001101010100110101010101010101010101000101001110101011111111101111111111111111111111111101111101011011010011111100001111111111111111111111111111111111111111111111111111111111111111111111111111111000111110011111101110110001,
	240'b101111001111111111001101010100110101010101010101010101010101001101010111101100001111111011111111111111111111101111000001101100001101011011111111111111111111111111111111111111111111111111111111111111111111111111111010111110111111101110110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010011010101111010010111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111110010110001,
	240'b101111001111111111001101010100110101010101010101010101010101010101010101010100110101001110001101111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111000011111111010110001,
	240'b101111001111111111001101010100110101010101010010010100100101010101010101010101010101010001010000011010101011010111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010010110110011111111110110001,
	240'b101111001111111111001101010100100101010110001110011111000101001001010101010101010101010101010101010100100101001101110110101100111110011011111110111111111111111111111111111111111111111111111111111110111010101001011010110111011111111110110001,
	240'b101111001111111111001101010100100101000010110010110100010101010101010100010101010101010101010101010101010101010101010001010100100110011010000111101011101100100111011001111000011110001011001100100011010101010001011001110111101111111110110001,
	240'b101111001111111111001101010100110101000101111001111011000111001001010010010101010101010101010101010101010101010101010101010101010101001101010001010100000101010001011101011000110110001101010111010100010101001101011010110111101111111110110001,
	240'b101111001111111111001101010100110101001101011000110110001010010101010000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010011010100110101001101010100010101010101010001011010110111101111111110110001,
	240'b101111001111111111001101010100110101001001001111101001001101100001011001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111001101010101010110001001010100011100001110101101111010010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101111001111111111001010011001101101100001110001010100001100110110110000010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111101111111110110001,
	240'b101110001111111111001100011010101111100111001011101101101110000111011011010110000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110111111111111110101101,
	240'b101000011111111111100100011101001100100011011001110110101101100110111000010110000101001101010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000100111101101111111100011111111010010100,
	240'b101001001111010011111111101110010110100001011101010111100101111001011101010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110010110100111000111111111111110110010011111,
	240'b110100011100100111111111111111111110010111010111110110001101100011011000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011110100111111111111111101100000111011000,
	240'b111100001100100011010001111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110001111100100111110001,
	240'b111101101111011111001001101011101011101011000100110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100010110000110100001111011111110110,
};
assign data = picture[addr];
endmodule