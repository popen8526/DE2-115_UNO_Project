module red_zero(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
    240'b111100101111101011100101101110101011000010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011000010110010110100011111000011101111,
    240'b111110101110011010111111111001101111110111111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011101110110000101100101011110010,
    240'b111010001100000011110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100010011010101,
    240'b101100111110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110111,
    240'b101000011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010,
    240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000,
    240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111,
    240'b101001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110,
    240'b101001101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111001,
    240'b110101101100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111000100,
    240'b111110001100111011010010111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011100111101011,
    240'b111110001111100111001000101110011100101011010001110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100011100110010111110101111001110110011110110,
    240'b111100111111101111100110101110111011000010110010101100101011001010110010101100101011001110110011101100111011001110110011101100101011001010110010101100101011001010110011101100111011001110110011101100111011000010110010110100101111000011101111,
    240'b111110101110011010111111111001101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110000101100100111110010,
    240'b111010001100000011110110111111111111111011110100111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111101011111111111111101100010011010101,
    240'b101100111110001011111111111000101000111101110100011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111000001101111011011101000000111001110111111111111010010110111,
    240'b101000011111101111111000100000000100110101010001010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010011110111000110100011100011100101010001100100111001011111111111000010,
    240'b101100101111111111011111010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011110011110110011101101111101111011001101010001101111001111111111000111,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101111101101100001100101100110011111000101101100101100101111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100011010111101001011011011001110101001111101101100101111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100011010111001001110011011101110100101111101101100101111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100101010110101001101011011001110100101111110101100101111111111001000,
    240'b101101101111111111011000010110100101010001010011010100000101001001010010010100000100111101010001010100110101010001010101010101010101010101010101010101010101010001010100110010001100011001010001100000011111000001110100101100101111111111001000,
    240'b101101101111111111011000010110100101000001100111100110101011000110110001101010011001011101111110011000110101010001010000010101000101010101010101010101010101010101010001100100001111011111001010111010011101000101010111101101011111111111000111,
    240'b101101101111111111011000010101111000010011100011111111111111111111111111111111111111111111111000111001011011111010001000010110110101000001010100010101010101010101010100010101111001100011010001101111000110101101001111101101101111111111000111,
    240'b101101101111111111010101011110111110110111111111111111111111111111111111111111111111111111111111111111111111111111111100110101001000110001010111010100100101010101010101010101000101001001010111010101000101001001010010101101101111111111000111,
    240'b101101101111111111011000110001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111000011011011010101000101010101010101010101010101010100010101000101010101010010101101101111111111000111,
    240'b101101101111111111101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111000011001010001010101000101010101010101010101010101010101010010101101101111111111000111,
    240'b101101101111111111110001111111001111111111111111111111111111111111111111111111111111111111111111111111111111110011101101111010101111100011111111111111111111010010010011010100010101010001010101010101010101010101010010101101101111111111000111,
    240'b101101101111111111110001111110111111111111111111111111111111111111111111111111111111111111111111110101001000100101100101011000100111110011000001111111001111111111110111100100010101000101010101010101010101010101010010101101101111111111001000,
    240'b101101101111111111110000111110111111111111111111111111111111111111111111111111111111111111000110010111110100111001001110010011100100111101010101101010001111110111111111111100111000000001010000010101010101010101010010101101101111111111001000,
    240'b101101101111111111101100111101101111111111111111111111111111111111111111111111111110100101101001010011110101100101111101100001000110000001010001010110001100110111111111111111111110001001101001010100100101010101010010101101101111111111001000,
    240'b101101101111111111100011111001111111111111111111111111111111111111111111111111111011000101001111010101101011000111111001111111101100110101100010010011011000110011111101111111111111111110111110010101010101010001010010101101101111111111001000,
    240'b101101101111111111011001110100111111111111111111111111111111111111111111111111111000101001001100011110101111100111111111111111111111111110011011010011010110110011110010111111111111111111111011100010000101000001010010101101101111111111001000,
    240'b101101101111111111010100101100111111111111111111111111111111111111111111111111100111110101001011100100001111111111111111111111111111111110110101010011110110010111101001111111111111111111111111110101010101101101010001101101101111111111000111,
    240'b101101101111111111010100100011101111110111111111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111011000101001001101101101101111111111000111,
    240'b101101101111111111010110011010101110011111111111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111100100101010010101101011111111111000111,
    240'b101101101111111111011000010110001011101111111111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111111001101101101101100111111111111000111,
    240'b101101101111111111011000010101100111111011111010111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111111111110011000101100011111111111000111,
    240'b101101101111111111011000010110010101011111001111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111111111111000010101101001111111111000111,
    240'b101101101111111111011000010110100100111110000011111110101111111111111111111111111000001001001011100001111111111111111111111111111111111110101011010011010110011111101110111111111111111111111111111111111111111111011111110000011111111111001000,
    240'b101101101111111111011000010110100101001101010101101111101111111111111111111111111001111001001101011000101101110011111111111111111111001001111000010011010111101111111010111111111111111111111111111111111111111111110001110100011111111111001000,
    240'b101101101111111111011000010110100101010001010010011010011110011011111111111111111101001001011001010100000111000110111001110000101000010001010011010100001011000011111111111111111111111111111111111111111111111111111010110111101111111111001000,
    240'b101101101111111111011000010110100101010001010101010100001000100011110101111111111111110010011100010100010101000001010011010101000101000001001111011111101111001011111111111111111111111111111111111111111111111111111100111001111111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101000110011101111110111111111111110111101000010101111001010001010100000101100010001001111010011111111111111111111111111111111111111111111111111111111111111100111011001111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010001010100101001001111101111111111111111111101110010110111101100111101000111111001111111111111111111111111111111111111111111111111111111111111111111111101111011111111111111000111,
    240'b101101101111111111011000010110100101010001010101010101010101010101010100010101001001101011110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001101111111111000111,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101000101000110000101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011101111111111000111,
    240'b101101101111111111011000010110100101010001010010010100000101001001010101010101010101010101010000011001011010111011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100101101011111111111000111,
    240'b101101101111111111011000010110100101001001110100100100110111010101010100010101010101010101010101010100100101001001110010101100001110010111111110111111111111111111111111111111111111111111111111111111111100111101100001101101001111111111000111,
    240'b101101101111111111011000010101111000011011110001111101011111001110001011010100010101010101010101010101010101010101010010010100100110010110001000101100001100111011011110111001111110101011011101101010010110000001001111101101101111111111000111,
    240'b101101101111111111010111010111101101011111000110011011011100001111011011010110110101010001010101010101010101010101010101010101010101001101010000010100010101010101100000011001110110101001011110010100010101001101010010101101101111111111001000,
    240'b101101101111111111010110011010001110011110001101010001111000100011101100011000110101001101010101010101010101010101010101010101010101010101010101010101010101010001010011010100110101001001010011010101010101010101010010101101101111111111001000,
    240'b101101101111111111010110011010011110011010001101010010111000011111101100011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101101111111111001000,
    240'b101101101111111111010110011010011110011010001100010010101000011011101100011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101101111111111001000,
    240'b101101101111111111010111011001001110011010011100010010011001100011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101101111111111001000,
    240'b101101011111111111011010010110001011100011101110101101011110110110111100010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101111111111111000111,
    240'b101001111111111111101110011001100101111110111011111000111011110101100100010100100101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001001010110110100101111111111000110,
    240'b101001101111000011111111101110100101111001010101010111100101011001010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011101111110101111110010111001,
    240'b110101101100100111111111111111111101111111001010110010011100101011001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010101101011011111011111111111101100111000100,
    240'b111110001100111011010010111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011100111101011,
    240'b111110001111100111001000101110011100101011010001110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100011100110010111110101111001110110011110110,
    240'b111100101111101011100101101110101011000010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011000010110010110100011111000011101111,
    240'b111110101110011010111111111001101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110000101100101011110010,
    240'b111010001100000011110110111111111111111011110100111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111101011111111111111101100010011010101,
    240'b101100111110001011111111111000101000111101110100011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111000001101111011011101000000111001110111111111111010010110111,
    240'b101000011111101111111000100000000100110101010001010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010011110111000110100011100011100101010001100100111001011111111111000010,
    240'b101100101111111111011111010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011110011110110011101101111101111011001101010001101111001111111111000111,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011101111101101100001100101100110011111000101101100101100101111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100011010111101001011011011001110101001111101101100101111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100011010111001001110011011101110100101111101101100101111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110110100101010110101001101011011001110100101111110101100101111111111001000,
    240'b101101101111111111011000010110100101010001010011010100000101001001010010010100000100111101010001010100110101010001010101010101010101010101010101010101010101010001010100110010001100011001010001100000011111000001110100101100101111111111001000,
    240'b101101101111111111011000010110100101000001100111100110101011000110110001101010011001011101111110011000110101010001010000010101000101010101010101010101010101010101010001100100001111011111001010111010011101000101010111101101011111111111000111,
    240'b101101101111111111011000010101111000010011100011111111111111111111111111111111111111111111111000111001011011111010001000010110110101000001010100010101010101010101010100010101111001100011010001101111000110101101001111101101101111111111000111,
    240'b101101101111111111010101011110111110110111111111111111111111111111111111111111111111111111111111111111111111111111111100110101001000110001010111010100100101010101010101010101000101001001010111010101000101001001010010101101101111111111000111,
    240'b101101101111111111011000110001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111000011011011010101000101010101010101010101010101010100010101000101010101010010101101101111111111000111,
    240'b101101101111111111101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111000011001010001010101000101010101010101010101010101010101010010101101101111111111000111,
    240'b101101101111111111110001111111001111111111111111111111111111111111111111111111111111111111111111111111111111110011101101111010101111100011111111111111111111010010010011010100010101010001010101010101010101010101010010101101101111111111000111,
    240'b101101101111111111110001111110111111111111111111111111111111111111111111111111111111111111111111110101001000100101100101011000100111110011000001111111001111111111110111100100010101000101010101010101010101010101010010101101101111111111001000,
    240'b101101101111111111110000111110111111111111111111111111111111111111111111111111111111111111000110010111110100111001001110010011100100111101010101101010001111110111111111111100111000000001010000010101010101010101010010101101101111111111001000,
    240'b101101101111111111101100111101101111111111111111111111111111111111111111111111111110100101101001010011110101100101111101100001000110000001010001010110001100110111111111111111111110001001101001010100100101010101010010101101101111111111001000,
    240'b101101101111111111100011111001111111111111111111111111111111111111111111111111111011000101001111010101101011000111111001111111101100110101100010010011011000110011111101111111111111111110111110010101010101010001010010101101101111111111001000,
    240'b101101101111111111011001110100111111111111111111111111111111111111111111111111111000101001001100011110101111100111111111111111111111111110011011010011010110110011110010111111111111111111111011100010000101000001010010101101101111111111001000,
    240'b101101101111111111010100101100111111111111111111111111111111111111111111111111100111110101001011100100001111111111111111111111111111111110110101010011110110010111101001111111111111111111111111110101010101101101010001101101101111111111000111,
    240'b101101101111111111010100100011101111110111111111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111011000101001001101101101101111111111000111,
    240'b101101101111111111010110011010101110011111111111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111100100101010010101101011111111111000111,
    240'b101101101111111111011000010110001011101111111111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111111001101101101101100111111111111000111,
    240'b101101101111111111011000010101100111111011111010111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111111111110011000101100011111111111000111,
    240'b101101101111111111011000010110010101011111001111111111111111111111111111111111010111110001001011100100011111111111111111111111111111111110110110010011110110010111101000111111111111111111111111111111111111111111000010101101001111111111000111,
    240'b101101101111111111011000010110100100111110000011111110101111111111111111111111111000001001001011100001111111111111111111111111111111111110101011010011010110011111101110111111111111111111111111111111111111111111011111110000011111111111001000,
    240'b101101101111111111011000010110100101001101010101101111101111111111111111111111111001111001001101011000101101110011111111111111111111001001111000010011010111101111111010111111111111111111111111111111111111111111110001110100011111111111001000,
    240'b101101101111111111011000010110100101010001010010011010011110011011111111111111111101001001011001010100000111000110111001110000101000010001010011010100001011000011111111111111111111111111111111111111111111111111111010110111101111111111001000,
    240'b101101101111111111011000010110100101010001010101010100001000100011110101111111111111110010011100010100010101000001010011010101000101000001001111011111101111001011111111111111111111111111111111111111111111111111111100111001111111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101000110011101111110111111111111110111101000010101111001010001010100000101100010001001111010011111111111111111111111111111111111111111111111111111111111111100111011001111111111001000,
    240'b101101101111111111011000010110100101010001010101010101010101010001010100101001001111101111111111111111111101110010110111101100111101000111111001111111111111111111111111111111111111111111111111111111111111111111111101111011111111111111000111,
    240'b101101101111111111011000010110100101010001010101010101010101010101010100010101001001101011110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001101111111111000111,
    240'b101101101111111111011000010110100101010001010101010101010101010101010101010101000101000110000101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011101111111111000111,
    240'b101101101111111111011000010110100101010001010010010100000101001001010101010101010101010101010000011001011010111011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100101101011111111111000111,
    240'b101101101111111111011000010110100101001001110100100100110111010101010100010101010101010101010101010100100101001001110010101100001110010111111110111111111111111111111111111111111111111111111111111111111100111101100001101101001111111111000111,
    240'b101101101111111111011000010101111000011011110001111101011111001110001011010100010101010101010101010101010101010101010010010100100110010110001000101100001100111011011110111001111110101011011101101010010110000001001111101101101111111111000111,
    240'b101101101111111111010111010111101101011111000110011011011100001111011011010110110101010001010101010101010101010101010101010101010101001101010000010100010101010101100000011001110110101001011110010100010101001101010010101101101111111111001000,
    240'b101101101111111111010110011010001110011110001101010001111000100011101100011000110101001101010101010101010101010101010101010101010101010101010101010101010101010001010011010100110101001001010011010101010101010101010010101101101111111111001000,
    240'b101101101111111111010110011010011110011010001101010010111000011111101100011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101101111111111001000,
    240'b101101101111111111010110011010011110011010001100010010101000011011101100011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101101111111111001000,
    240'b101101101111111111010111011001001110011010011100010010011001100011101001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101101111111111001000,
    240'b101101011111111111011010010110001011100011101110101101011110110110111100010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101111111111111000111,
    240'b101001111111111111101110011001100101111110111011111000111011110101100100010100100101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001001010110110100101111111111000110,
    240'b101001101111000011111111101110100101111001010101010111100101011001010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011101111110101111110010111001,
    240'b110101101100100111111111111111111101111111001010110010011100101011001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010101101011011111011111111111101100111000100,
    240'b111110001100111011010010111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011100111101011,
    240'b111110001111100111001000101110011100101011010001110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100011100110010111110101111001110110011110110,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule