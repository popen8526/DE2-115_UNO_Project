module red_nine(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111100001111001111110011110011101011010110110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011010111001000111010111111001011110000,
	240'b111100011110101011000010110100011111000011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111000111010010101110011110010011110001,
	240'b111011011011110111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011101111101100,
	240'b101110001100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010010111001,
	240'b100101101110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110010100,
	240'b101010111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010101001,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111,
	240'b101100101111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110001,
	240'b100111001111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110011010,
	240'b101000111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110100011,
	240'b110111111011101111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011111011011110,
	240'b111100101101011111000000111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110000001101000111110010,
	240'b111101111111101011011101101010011010011110111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010100010101001110110111111101011110111,
	240'b111100001111001111110100110011111011011010110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011010111001000111011001111001011110000,
	240'b111100011110101011000010110100011111000011110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111000111010010101110001110010011110001,
	240'b111011011011110111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011101111101100,
	240'b101110001100111011111111111101011011001010001101100010111000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000100110000111100010101010110111110010111111111101010010111001,
	240'b100101101110111011111110101000000100111101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010011100110100110000111011010010100110010010101111111011111011110010100,
	240'b101010111111110011110000011001110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000001110101111110101111011000111111001011110111001111111111110101001,
	240'b101110001111111111101000011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100101100101101110100110010111101000101100000110111101111111110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100001111001011001010101000001100101001110001101101000110111011111111110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111001101101011010001010110110011100100001011110110111101111111110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111000111111001111110010110110110111001001011010110111111111111110110111,
	240'b101110001111111111101000011000100101001101010100010100000101000001010001010100000101000001010010010101000101010101010101010101010101010101010101010101010101001101011110111000011010101101110001011101000101100101011101110111111111111110110111,
	240'b101110001111111111101000011000100101000001011100100001101001111010011110100101101000010101110000010110100101000101010001010101000101010101010101010101010101010101010010101101101110110110110001111001001001010101011001110111111111111110110111,
	240'b101110001111111111101000010111110110111111010000111111001111111111111111111111111111110111110000110101101010101001110110010101000101000101010101010101010101010101010011011000111011101011100000101110100110001101011100110111111111111110110111,
	240'b101110001111111111100101011100101101101111111111111111111111111111111111111111111111111111111111111111111111111111110011110000000111100001010010010100110101010101010101010100110101010101011110010101010101000101011101110111111111111110110111,
	240'b101110001111111111100100101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101010010111100101000101010101010101010101010001010011010101000101001101011101110111111111111110110111,
	240'b101110001111111111101111111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100110111101010000010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111110110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011110011111100101111110111111111111111111110001101111001010100000101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111110110111110111111111111111111111111111111111111111111111111111111111111111111110110011000111101101011011010101000101111010011111111111111111111100110011101010101000101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111110101111110111111111111111111111111111111111111111111111111111111111111001001011000010100111001001110010011100100111001011101110000001111111111111111110111100110100001010010010101010101001101011101110111111111111110110111,
	240'b101110001111111111110010111100101111111111111111111111111111111111111111111111111110101001101011010011110101100001111001011110110101101001001111011001001110001011111111111111111100010101011000010101000101001101011101110111111111111110110111,
	240'b101110001111111111101100111000001111111111111111111111111111111111111111111111111011001001001111010101111011001111111001111110101011110001011010010011101010011011111111111111111111111010011010010100000101001101011101110111111111111110110111,
	240'b101110001111111111100101110010111111111111111111111111111111111111111111111111111000101101001100011111101111101111111111111111111111111110000111010010111000000011111100111111111111111111101010011010110101000001011101110111111111111110110111,
	240'b101110001111111111100010101010101111111111111111111111111111111111111111111111100111110101001011100101011111111111111111111111111111111110011111010011000111100011110111111111111111111111111111101100010101000001011101110111111111111110110111,
	240'b101110001111111111100100100001111111100011111111111111111111111111111111111111010111110001001101011111001111101011111111111111111111111010000101010010111000001011111101111111111111111111111111111011100110100101011010110111111111111110110111,
	240'b101110001111111111100110011010101101101111111111111111111111111111111111111111010111110001010000010101101010101111110101111101111011010001011000010011101010101011111111111111111111111111111111111111111010000101011000110111111111111110110111,
	240'b101110001111111111101000010111101010101111111111111111111111111111111111111111010111110001010001010101000101011001110011011101010101011101001111011010011110011111111111111111111111111111111111111111111101011001100010110111101111111110110111,
	240'b101110001111111111101000010111100111001011110101111111111111111111111111111111010111110001010001010101010101000001001110010011100100111001100010110010011111111111111111111111111111111111111111111111111111011001111111110110111111111110110111,
	240'b101110001111111111101000011000010101001011000010111111111111111111111111111111010111110001001101100000011001100101110011011100101001001011011001111111111111111111111111111111111111111111111111111111111111111110100011110110011111111110110111,
	240'b101110001111111111101000011000100100111101111000111101011111111111111111111111111000001101001011100011111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110110111011111111110110111,
	240'b101110001111111111101000011000100101001101010011101100101111111111111111111111111001111101001101011001001101111011111111111111111110000110011110110111101111110111111111111111111111111111111111111111111111111111100001111000011111111110110111,
	240'b101110001111111111101000011000100101001101010010011000101101110111111111111111111101010101011001010100000111000110110101101101100111010001001101011001101110001011111111111111111111111111111111111111111111111111101101111010011111111010110111,
	240'b101110001111111111101000011000100101001101010101010100010111110111110001111111111111110110011111010100010101000001010010010100100101000001001111100100001111100011111111111111111111111111111111111111111111111111110011111100011111110110110111,
	240'b101110001111111111101000011000100101001101010101010101010101000010010011111110001111111111110111101001100110010101010101010101010110000010011011111100111111111111111111111111111111111111111111111111111111111111110110111101001111110110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010001010001100110011111100011111111111101011100010010100100101000011100000011110001111111111111111111111111111111111111111111111111111111111111111111110111111101101111110010110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010100010100101001000111110010110011000111001101110110011101100111001010111111111111111111111111111111111111111111111111111111111111111111111111110010111011101111110110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101000101000101111101110011101110101011101010111010001110011111110100111111111111111111111111111111111111111111111111111111111111111111010110111000001111111110110111,
	240'b101110001111111111101000011000100101001101010001010100010101000101010100010101010101010101010000011000011010011111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001111110110111111111110110111,
	240'b101110001111111111101000011000100101001001111011101000111000011001010110010101000101010101010101010100110101000101101011101001011101110111111010111111111111111111111111111111111111111111111111111110001010001001011100110111101111111110110111,
	240'b101110001111111111101000010111101000001011110011111011001111011110011010010100100101010101010101010101010101010101010010010100010101111101111100101000111011111111010001110110101101101111000100100001010101001001011100110111111111111110110111,
	240'b101110001111111111101000011000000110110110010101011001001010110111100011010111010101001101010101010101010101010101010101010101010101001101010001010100000101001001011001010111100101111001010101010100010101001001011101110111111111111110110111,
	240'b101110001111111111101000011000010101010110011101110010011100101011101110011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010100010100110101001101010100010101010101001101011101110111111111111110110111,
	240'b101110001111111111101000010111101001110111110101110011101111001011110000011000110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111100111011001001101100110101111010010111001011111110001011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111100111011000111101011110110011010011111001110011101001010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101100101111111111101011010111111001100111110110110100011111001110110000010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111000011111111110110001,
	240'b100111001111010111111010011111110101000010011000110010101010010001011011010100100101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110100111001110111111101011111110110011010,
	240'b101000111101111011111111110110010111011101011101011000000101110101011111011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000000111010011010010111111111110010110100011,
	240'b110111111011101111111000111111111111010011100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011111001011111111111110101011111011011110,
	240'b111100101101011111000000111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110000001101000111110010,
	240'b111101111111101011011101101010011010011110111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010100010101001110110111111101011110111,
	240'b111100001111001111110011110011101011010110110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011010111001000111010111111001011110000,
	240'b111100011110101011000010110100011111000011110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111000111010010101110011110010011110001,
	240'b111011011011110111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011101111101100,
	240'b101110001100111011111111111101011011001010001101100010111000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000100110000111100010101010110111110010111111111101010010111001,
	240'b100101101110111011111110101000000100111101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010011100110100110000111011010010100110010010101111111011111011110010100,
	240'b101010111111110011110000011001110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000001110101111110101111011000111111001011110111001111111111110101001,
	240'b101110001111111111101000011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010111110100101100101101110100110010111101000101100000110111101111111110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100001111001011001010101000001100101001110001101101000110111011111111110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111001101101011010001010110110011100100001011110110111101111111110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100010111000111111001111110010110110110111001001011010110111111111111110110111,
	240'b101110001111111111101000011000100101001101010100010100000101000001010001010100000101000001010010010101000101010101010101010101010101010101010101010101010101001101011110111000011010101101110001011101000101100101011101110111111111111110110111,
	240'b101110001111111111101000011000100101000001011100100001101001111010011110100101101000010101110000010110100101000101010001010101000101010101010101010101010101010101010010101101101110110110110001111001001001010101011001110111111111111110110111,
	240'b101110001111111111101000010111110110111111010000111111001111111111111111111111111111110111110000110101101010101001110110010101000101000101010101010101010101010101010011011000111011101011100000101110100110001101011100110111111111111110110111,
	240'b101110001111111111100101011100101101101111111111111111111111111111111111111111111111111111111111111111111111111111110011110000000111100001010010010100110101010101010101010100110101010101011110010101010101000101011101110111111111111110110111,
	240'b101110001111111111100100101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101010010111100101000101010101010101010101010001010011010101000101001101011101110111111111111110110111,
	240'b101110001111111111101111111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100110111101010000010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111110110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011110011111100101111110111111111111111111110001101111001010100000101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111110110111110111111111111111111111111111111111111111111111111111111111111111111110110011000111101101011011010101000101111010011111111111111111111100110011101010101000101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111110101111110111111111111111111111111111111111111111111111111111111111111001001011000010100111001001110010011100100111001011101110000001111111111111111110111100110100001010010010101010101001101011101110111111111111110110111,
	240'b101110001111111111110010111100101111111111111111111111111111111111111111111111111110101001101011010011110101100001111001011110110101101001001111011001001110001011111111111111111100010101011000010101000101001101011101110111111111111110110111,
	240'b101110001111111111101100111000001111111111111111111111111111111111111111111111111011001001001111010101111011001111111001111110101011110001011010010011101010011011111111111111111111111010011010010100000101001101011101110111111111111110110111,
	240'b101110001111111111100101110010111111111111111111111111111111111111111111111111111000101101001100011111101111101111111111111111111111111110000111010010111000000011111100111111111111111111101010011010110101000001011101110111111111111110110111,
	240'b101110001111111111100010101010101111111111111111111111111111111111111111111111100111110101001011100101011111111111111111111111111111111110011111010011000111100011110111111111111111111111111111101100010101000001011101110111111111111110110111,
	240'b101110001111111111100100100001111111100011111111111111111111111111111111111111010111110001001101011111001111101011111111111111111111111010000101010010111000001011111101111111111111111111111111111011100110100101011010110111111111111110110111,
	240'b101110001111111111100110011010101101101111111111111111111111111111111111111111010111110001010000010101101010101111110101111101111011010001011000010011101010101011111111111111111111111111111111111111111010000101011000110111111111111110110111,
	240'b101110001111111111101000010111101010101111111111111111111111111111111111111111010111110001010001010101000101011001110011011101010101011101001111011010011110011111111111111111111111111111111111111111111101011001100010110111101111111110110111,
	240'b101110001111111111101000010111100111001011110101111111111111111111111111111111010111110001010001010101010101000001001110010011100100111001100010110010011111111111111111111111111111111111111111111111111111011001111111110110111111111110110111,
	240'b101110001111111111101000011000010101001011000010111111111111111111111111111111010111110001001101100000011001100101110011011100101001001011011001111111111111111111111111111111111111111111111111111111111111111110100011110110011111111110110111,
	240'b101110001111111111101000011000100100111101111000111101011111111111111111111111111000001101001011100011111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110110111011111111110110111,
	240'b101110001111111111101000011000100101001101010011101100101111111111111111111111111001111101001101011001001101111011111111111111111110000110011110110111101111110111111111111111111111111111111111111111111111111111100001111000011111111110110111,
	240'b101110001111111111101000011000100101001101010010011000101101110111111111111111111101010101011001010100000111000110110101101101100111010001001101011001101110001011111111111111111111111111111111111111111111111111101101111010011111111010110111,
	240'b101110001111111111101000011000100101001101010101010100010111110111110001111111111111110110011111010100010101000001010010010100100101000001001111100100001111100011111111111111111111111111111111111111111111111111110011111100011111110110110111,
	240'b101110001111111111101000011000100101001101010101010101010101000010010011111110001111111111110111101001100110010101010101010101010110000010011011111100111111111111111111111111111111111111111111111111111111111111110110111101001111110110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010001010001100110011111100011111111111101011100010010100100101000011100000011110001111111111111111111111111111111111111111111111111111111111111111111110111111101101111110010110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010100010100101001000111110010110011000111001101110110011101100111001010111111111111111111111111111111111111111111111111111111111111111111111111110010111011101111110110110111,
	240'b101110001111111111101000011000100101001101010101010101010101010101010101010101000101000101111101110011101110101011101010111010001110011111110100111111111111111111111111111111111111111111111111111111111111111111010110111000001111111110110111,
	240'b101110001111111111101000011000100101001101010001010100010101000101010100010101010101010101010000011000011010011111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001111110110111111111110110111,
	240'b101110001111111111101000011000100101001001111011101000111000011001010110010101000101010101010101010100110101000101101011101001011101110111111010111111111111111111111111111111111111111111111111111110001010001001011100110111101111111110110111,
	240'b101110001111111111101000010111101000001011110011111011001111011110011010010100100101010101010101010101010101010101010010010100010101111101111100101000111011111111010001110110101101101111000100100001010101001001011100110111111111111110110111,
	240'b101110001111111111101000011000000110110110010101011001001010110111100011010111010101001101010101010101010101010101010101010101010101001101010001010100000101001001011001010111100101111001010101010100010101001001011101110111111111111110110111,
	240'b101110001111111111101000011000010101010110011101110010011100101011101110011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010100010100110101001101010100010101010101001101011101110111111111111110110111,
	240'b101110001111111111101000010111101001110111110101110011101111001011110000011000110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111100111011001001101100110101111010010111001011111110001011001000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101110001111111111100111011000111101011110110011010011111001110011101001010111110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110111,
	240'b101100101111111111101011010111111001100111110110110100011111001110110000010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111000011111111110110001,
	240'b100111001111010111111010011111110101000010011000110010101010010001011011010100100101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110100111001110111111101011111110110011010,
	240'b101000111101111011111111110110010111011101011101011000000101110101011111011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000000111010011010010111111111110010110100011,
	240'b110111111011101111111000111111111111010011100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011111001011111111111110101011111011011110,
	240'b111100101101011111000000111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110000001101000111110010,
	240'b111101111111101011011101101010011010011110111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010100010101001110110111111101011110111,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule