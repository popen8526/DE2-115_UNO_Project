module Uno();
// None, because this is a top module.
endmodule