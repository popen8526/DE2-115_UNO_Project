module Player();
endmodule