module yellow_draw_two(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110101111110011100101100110011001010110110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100001000111110101001111100101111110011111010,
	240'b111111111111100010111111110010101101110111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000101101101111000111110011011111110111111111,
	240'b111111101100010011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001100111011111111,
	240'b110011101101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100011001101,
	240'b101000011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110011111,
	240'b101010111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110000,
	240'b101100011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111100011011010110110011101101011011010110110011101110111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111100011111001101110110011101100111011001110110011101011011001001111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111100100011110101111111111111111111111111111111111111111111010110111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111101101011011110111111111111111111111111111111111111111111101010110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111110110011001110111111111111111111111111111111111111111111111011101110011101100011011010111001001111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111101011000110111111011111111111111111111111111111111111111111101111101100100111011000110011101101001011111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111001100111011111111111111111111111111111111111111111111110110101110010011111111111111111100101011101111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111011011110111101111111111111111111111111111111111111111111011011100111011111111111111111101101111011101111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111101101110011011111111111111111111111111111111111111111111110011100011111111100111111111110111111001011111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111011110001101111110011111111111111111111111111111111111111111100101011110001111111111111101111000111111110101111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111110011001110111111111111111111111111111111111111111111111101101111011110111111111111111111001100111011111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111110110111101110011111111111111111111111111111111111111111110111011001111111111111111111111011110110110111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111101001100011011100011111001111110011111100111111010001101100111000100111111111111111111101111110011011111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111110111011010001110011111100100010101010110100001100110111101101111111111111111111111100110001011111101111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001000111110111111111111111111111111111111111111111111110011101110110011111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001101111011011111111111111111111111111111111111111111111000001101101111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001110010011110110011101111111011111110111111110000110110001100101111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100101011001001110010011100100111001001110010011111001011111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101100101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110110,
	240'b101011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110100,
	240'b101000011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010100010,
	240'b101110001101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000110110101,
	240'b111101011011111111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101100001111110111,
	240'b111111101110011010111100111001101111110111111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011011110101111011111000011111110,
	240'b111100011111010011101000101011011010011010101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011101010010010101111111010001111001111110001,
	240'b111110101111110011100101100110011001010110110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100001000111110101001111100101111110011111010,
	240'b111111111111100010111111110010101101110111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000101101101111000111110011011111110111111111,
	240'b111111101100010011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001100111011111111,
	240'b110011101101001011111111111110111101110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011101100110111001110110011111100111111001111110100001110001111111110111111111100100011001101,
	240'b101000011111010011111110110011101010100010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100110101011001011101110110100101001101010011110100111101001111010101011011010111111111110010110011111,
	240'b101010111111111111110100101100011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111001111111101111110110110010001010100010101010101010101010011110111010111111001111010110110000,
	240'b101100011111111111101110101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011010100111101001100001011011100111101011011000110101001101010001010011110110110111110001111011110110110,
	240'b101100101111111111101110101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011100100110111011010010010110100111001001011010110101001110011101011010010110011111110001111011110110110,
	240'b101100101111111111101110101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011010100111100111011011010100111101010111010110110111111111110001101000010111100111110001111011110110110,
	240'b101100101111111111101110101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111001101111001110111111101001101011100011110111111111111111101111011011111101011111011110110110,
	240'b101100101111111111101110101011101010100110101001101010001010011110101000101010001010100010101001101010101010101010101010101010101010101010101110101100101101110011110111110100001010111111000101111110011101010110111111111101111111011110110110,
	240'b101100101111111111101110101011101010011110101101110000011100110011001011110001111011110010110010101010101010100010101001101010101010100011100000111001101101000111110100111111111011100110101010110101001011011010110011111110001111011110110110,
	240'b101100101111111111101110101011001011100011101000111111011111111111111111111111111111110011110011111000111100101110110100101010001010011111011010111100111111000111110000111011101011011110101000101010011010100010110110111110001111011110110110,
	240'b101100101111111111101101101110001111000011111111111111111111111111111111111111111111111111111111111111111111111111110100110101111011010010101100101100001011000110110001101100001010101110101010101010101010100010110110111110001111011110110110,
	240'b101100101111111111101101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111001010101010101010100010101001101010011010101010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111011110011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101011000010101000101010101010101010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111011111000111110111111111111111111111111111111100011011010110110011101101011011010110110011101110111111001111111111111111111111111111111111110100010110100101010001010101010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111011111001111111001111111111111111111111111100011111001101110110101101100111011001110110101101011111001001111110101111111111111111111111111111111111101011101100111010100010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111011110111111110111111111111111111111111111100100111110101111001101100110111001101110100001111000011010111111000001111111111111111111111111111111111111111111001101010111010101001101010101010100010110110111110001111011110110110,
	240'b101100101111111011110101111110011111111111111111111111111101101111011101110000101010010110101000101001101011100111100010110100101111111111111111111111111111111111111111111111111101100010101001101010101010100010110110111110001111011110110110,
	240'b101100101111111011110001111101001111111111111111111111111110110011010000110100011010011110101010101010101010101111100011101111001101100111011010111001001111111111111111111111111111110011000010101010001010100010110110111110001111011110110110,
	240'b101100101111111111101110111010011111111111111111111111111111101011001000111000001010101010101010101010101010011111010111110000011100101011011011110011111101001011111111111111111111111111101101101011111010100010110110111110001111011110110110,
	240'b101100101111111111101011110110011111111111111111111111111111111111001110111000111011001010101001101010101010100011000101110101101011110111011011111101111100101111101111111111111111111111111111110011011010011010110110111110001111011110110110,
	240'b101100101111111111101100110001101111111011111111111111111111111111011011110111001100000110101000101010101010100110110101111000111001011010100110110010001101101011011110111111111111111111111111111011111010110110110101111110001111011110110110,
	240'b101100101111111111101101101101011111001011111111111111111111111111101101110011111101001110100111101010101010101010101011111000111010010110100101101100111110010011001101111111111111111111111111111111101100010010110011111110001111011110110110,
	240'b101100101111111111101110101011001101101111111111111111111111111111111011110010011101111110101010101010101010101010101000110110001011101010011111101010111110000011001001111110101111111111111111111111111101111110110101111110001111011110110110,
	240'b101100101111111111101110101011001011110111111100111111111111111111111111110011011110010010110011101001111010100010100110110001001101010110011000101010011101001111001110111011111111111111111111111111111111001110111110111101111111011110110110,
	240'b101100101111111111101110101011101010101011100101111111111111111111111111110111001101110111100010101111011011110010111011110110001110111110011001101010001100000111011100110110111111111111111111111111111111110111001110111101011111011110110110,
	240'b101100101111111111101110101011101010011110111111111111001111111111111111111101001100011111100100111001001110001111100100111001111101101110010101101010001011001011100011110011101111111111111111111111111111111111011110111101011111011110110110,
	240'b101100101111111111101110101011101010100110101001110111001111111111111111111111111110111011010001110100001100100010101101101101111001001010100000101010111010101011011111110010001111101111111111111111111111111111101100111101111111011110110110,
	240'b101100101111111111101110101011101010100110101001101100101111000111111111111111111111111111111111111111111111110111001010111000101010101110101001101010001010010111010010110100001110110011111111111111111111111111110101111110001111011010110110,
	240'b101100101111111111101110101011101010100110101010101010001100000111111001111111111111111111111111111111111111111111001110111010101101000110110110101101101011010111011111111000101101101111111111111111111111111111111001111110101111011010110110,
	240'b101100101111111111101110101011101010100110101010101010101010100011001100111111001111111111111111111111111111111111101001110010101110110011101010111010101110101011101111110110001100101111111111111111111111111111111010111110111111011010110110,
	240'b101100101111111111101110101011101010100110101010101010101010101010101001110011101111110011111111111111111111111111111111111000111100101111001001110010101100101011001001110010011111001011111111111111111111111111111010111110111111011010110110,
	240'b101100101111111111101110101011101010100110101010101010101010101010101001101010011100100111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110011111011010110110,
	240'b101100101111111111101110101011101010100110101010101010101010101010101010101010011010100010111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010111101101111011110110110,
	240'b101100101111111111101110101011101010100110101010101010101010100110101000101010001010100010100110101011011100110111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011000001111101101111011110110110,
	240'b101100101111111111101110101011101010100010101000101010011011110011011111110111111110000111100000110000111010011010110010110010111110100011111001111111111111111111111111111111111111111111111111111100111011111110110100111110001111011110110110,
	240'b101100101111111111101110101011011011010010111100101001111100100011111111111100101110011011111010110101101010011110101001101010001010110010111001110010011101011111100001111001011110010011010100101101101010011110110110111110001111011110110110,
	240'b101100101111111111101110101011111101010111101010101011101011011111101110111100111100001010111100101110001010100110101010101010101010100110101000101010001010100010101001101010111010101010101000101010011010100010110110111110001111011110110110,
	240'b101100101111111111101101110110111111100111111101111010001010111010110000111000001111100111000110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111111101110110001111110101011110110110011111010110110100110101010111101010011111000101111001010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111111101110101010111100011111011011101001111011011111001010101010101010101011101101110101001010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110110111110001111011110110110,
	240'b101100101111111111101110101011101010101110101101101010001100000111111010101111101011010111110011110011111010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110110111110001111011110110110,
	240'b101011111111111111110001101011111010100110101001101010011010110111100101111110011111011011101111101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110111111110101111011110110100,
	240'b101000011111100111111100101111111010011010101000101010001010011110110000110011101101000110110100101001111010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011011001100111111111110110010100010,
	240'b101110001101111011111111111100001100010110111010101110101011101010111001101110001011100010111001101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100101111110111111111111101000110110101,
	240'b111101011011111111110100111111111111111011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111010101100001111110111,
	240'b111111101110011010111100111001101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011011110101111011111000011111110,
	240'b111100011111010011101000101011011010011010101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011101010010010101111111010001111001111110001,
	240'b111110101111110011100101100110011001010110110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101100001000111110101001111100101111110011111010,
	240'b111111111111100010111111110010101101110111100011111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111000101101101111000111110011011111110111111111,
	240'b111111101100010011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001100111011111111,
	240'b110011101101001011111111111100111001100101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011010110100101101011011011110110111101101111011100101010101011111011111111111100100011001101,
	240'b101000011111010011111101011011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011001000011101000000000000000000000000000000000000010010010001111111111110011010011111,
	240'b101010111111111111011101000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000101101101111001011100101010110100000000000000000000000000000000000110000111101001111011110110000,
	240'b101100011111111111001011000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110110111100100101110010101111000100001011100000000000000000000000000100010111010001111100110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101111100110110000000000011101101011010010000100000001011011010001111100011100111010001111100110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110110110100010010100000000000000110000101001000000111010100111001000110110111001111111100110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010101101001101100101000001000000000010100111100111111111101111001110010011111000011111100110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000110101001011111100111011100110001000101010000111011011000000000111111111001101111100110110110,
	240'b101100101111111111001011000011000000000000001011010001000110011001100100010101100011010100011001000000000000000000000000000000000000000010100000101101000111010011011111111111110010110000000000011111100010010100011100111010001111100110110110,
	240'b101100101111111111001011000001110010110110111010111110101111111111111111111111101111011111011011101010110110010000011101000000000000000010010000110110111101011011010011110011000010100100000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111000111001010111101000111111111111111111111111111111111111111111111111111111111111111111111111111011111100001110010000000001000000101000001010100010100000100110000010000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111000111100110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001100000000000010000000000000000000000000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111011010111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100111010001010100000000000000000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111101001111101001111111111111111111111111111100011011010110110101101101011011011110110101101110111111001111111111111111111111111111111111011101000011111000000000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111101011111101011111111111111111111111111100011111001101110111011101101011011010110110111101101111001010111110101111111111111111111111111111111111000010000111000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111100111111100101111111111111111111111111100100111110110101010100110001101100011011011001100011011011010111000001111111111111111111111111111111111111111101101000000111000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111100000111011111111111111111111111111111101110011011010010000110000000000000000000000000010100011010100110101001111111111111111111111111111111111111111111111111000100100000001000000000000000000100011111010001111100110110110,
	240'b101100101111111111010110110111011111111111111111111111111110110011010100011100000000000000000000000000000000000110110011110000001101100111011010111001001111111111111111111111111111011001001000000000000000000000100011111010001111100110110110,
	240'b101100101111111111001100101111001111111111111111111111111111101111001101101001110000000000000000000000000000000010000001110001011100110011011111110100011101001011111111111111111111111111001000000011110000000000100011111010001111100110110110,
	240'b101100101111111111000011100010111111111111111111111111111111111111010001110010010001010100000000000000000000000001001011110011110110111110000110111000011100110111101111111111111111111111111111011010010000000000100011111010001111100110110110,
	240'b101100101111111111000100010101001111101111111111111111111111111111011100110110000011111000000000000000000000000000011101110100000010100000000000010100111101100111011110111111111111111111111111110011110000101100100000111010001111100110110110,
	240'b101100101111111111001000001000001101100011111111111111111111111111101101110100110111010100000000000000000000000000000011101101110110001000000000000101101100110011010000111111111111111111111111111111010100111000011011111010001111100110110110,
	240'b101100101111111111001011000001111001001111111111111111111111111111111011110011101010011100000001000000000000000000000000100001001001101100000000000000011010100111001111111110101111111111111111111111111010000000100000111001111111100110110110,
	240'b101100101111111111001011000001010011100111110110111111111111111111111111110100001100111000010110000000000000000000000000010010001100100100001100000000000111010111010011111011111111111111111111111111111101110100111101111001001111100110110110,
	240'b101100101111111111001011000010100000010010110001111111111111111111111111110111001101110110011011001101100011000100110000011111111111000100101110000000000100000011010111110111001111111111111111111111111111100001101011111000011111100110110110,
	240'b101100101111111111001011000011000000000000111111111101011111111111111111111101001100011111100101110111101101110011011100111001011101111000111001000000000001010111001010110100011111111111111111111111111111111110011100111000011111100110110110,
	240'b101100101111111111001011000011000000000000000010100101101111111111111111111111111110111011010001110100011100101010110001100001010010000000000100000000000000000110100110110011011111101111111111111111111111111111000110111001011111100010110110,
	240'b101100101111111111001011000011000000000000000000000110101101010011111111111111111111111111111111111111111111110111001111101100010000000000000000000000000000000001110010110101001110110011111111111111111111111111100011111010011111100010110110,
	240'b101100101111111111001011000011000000000000000000000000000100010111101110111111111111111111111111111111111111111111001111111000110110111100100011001000100010001110010101111001001101101111111111111111111111111111101101111011101111011110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000001100110111101111111111111111111111111111111111111101000110010111110101111100000110111111110000011101101110110001100101111111111111111111111111111101111111100011111011110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000011011011111011011111111111111111111111111111111111000111100101111001011110010111100101111001001110010011111001011111111111111111111111111110001111100011111011110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000101110111101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111010111111100010110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000000000000110111101110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001111000101111100110110110,
	240'b101100101111111111001011000011000000000000000000000000000000000000000000000000000000000000000000000010100110101011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101000110111000111111100110110110,
	240'b101100101111111111001011000011000000000000000000000000000011010110011110101000011010010010100011010011010000000000011010011001011011101111101110111111111111111111111111111111111111111111111111110110110100000000011101111010001111100110110110,
	240'b101100101111111111001011000010000010000100110111000000000101101111111111110110011011010011110001100001000000000000000000000000000000011100101101010111011000100010100100101100001010111101111111001001000000000000100011111010001111100110110110,
	240'b101100101111111111001011000100001000000011000001000011110010100011001011110110110100011000110101001010100000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111001001100101001110110111111000101110110000110000010110101000101110110001010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111001010010110001011111111100101011011010000011100000000000001010111110111101010001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111001011000000110101100110010010000000000010100001100000000000000000000011001010011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111010001111100110110110,
	240'b101100101111111111001010000010110000010100001000000000000100010111110001001110110010000011011011011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111010001111100110110110,
	240'b101011111111111111010011000011100000000000000000000000000000110010110011111011001110010011010001000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110111011101111100110110100,
	240'b101000011111101011110101010000000000000000000000000000000000000000010001011010110111011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101111111101110110010100010,
	240'b101110001101111011111111110100100101000100101111001100000011000000101101001010100010101000101100001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100010110001011100101111111111101000110110101,
	240'b111101011011111111110100111111111111110011101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101111111111111111111010101100001111110111,
	240'b111111101110011010111100111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011110101111011111000011111110,
	240'b111100011111010011101000101011011010011010101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011101010010010101111111010001111001111110001,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule