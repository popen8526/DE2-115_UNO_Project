module blue_six(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111111111111101011100100101000001001101010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101011111001011110110100111110111111111111111111,
	240'b111111111110110010110110110101101111010111110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111001011001111110001001111100111111111,
	240'b111110111100000111100111111111111111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111111111111111111111110111001100110011111011,
	240'b110001101101011011111111111100001010100110001010100010011000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010011000011010000101100010101011010011111000111111111100110011000010,
	240'b100011111111010011111101100101100100111001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010100010111010110001011011000110100111010101110111111111110001110010101,
	240'b101000011111110011101011011000110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100110011111010111110100111000100110101101110010111110111110111110100010,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100100001001111001110011110111001011010101101000111101111111010110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010110101001100110101101110100011100110101101010111101111111010110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100101100101111011011100011111111111100101101101010111101111111010110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100110111011101001010101011001110010101101000001101010111101111111010110110000,
	240'b101100011111111111100100010111010101001101010011010100000101000001010000010011110101000001010010010101000101010101010101010101010101010101010101010101010101001001101011111100011000000101001001101110111100101001101010111101111111010110110000,
	240'b101100011111111111100100010111010100111101100000100010101010001010100001100101011000001101101100010110000101000001010010010101000101010101010101010101010101010001011000110010111110010010111011111101011001010101101000111101111111010110110000,
	240'b101100011111111111100100010110010111100011011000111111101111111111111111111111111111101111101110110100101010010101110010010100110101000101010101010101010101010101010010011011001100010111100000101001110101011001101011111101111111010110110000,
	240'b101100011111111111100010011100101110001111111111111111111111111111111111111111111111111111111111111111111111111111110001101110100111000101010001010101000101010101010101010100100101011001011101010100110101000101101100111101111111010110110000,
	240'b101100011111111111100000101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110100000010110000101001001010101010101010101010001010011010101010101001001101100111101111111010110110000,
	240'b101100011111110111101101111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000100110001101010001010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100011111110011111010111101111111111111111111111111111111111111111111111111111111111111111111111111111111110011110010111100111111111011111111111111111101010001101010010100010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100011111110011111011111110011111111111111111111111111111111111111111111111111111111111111111110011101000011101101001011010111001000011011100111111111111111111011000011010000101001001010101010101010101001001101100111101111111010110110000,
	240'b101100011111110011111000111101011111111111111111111111111111111111111111111111111111111110111011010110110100111101001110010011100100111001100101110100001111111111111111110011010101110001010011010101010101001001101100111101111111010110110000,
	240'b101100011111110111110011111011101111111111111111111111111111111111111111111111111110001001011111010011100101101001111100011110010101011101001110011100011111000011111111111111111010111001010011010101010101001001101100111101111111010110110000,
	240'b101100011111111011101001111000011111111111111111111111111111111111111111111111111111000110100100011010011011110011111011111110001010110001010101010100011011110111111111111111111111100010000011010100000101001001101100111101111111010110110000,
	240'b101100011111111011100010110011011111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111110001110111010011001001011111111111111111111111111111011000010111000101000001101100111101111111010110110000,
	240'b101100011111111111011111101010111111111111111111111111111111111111111111111111111111111111111111111111001100111010101101101011101101011010001010010011001000101011111111111111111111111111111111100101100100110101101100111101111111010110110000,
	240'b101100011111111111100000100010011111101011111111111111111111111111111111111111111111111111101011100010100101011101010000010100000101110001011111010011111000100111111111111111111111111111111111110110100101100101101011111101111111010110110000,
	240'b101100011111111111100011011010001110001011111111111111111111111111111111111111111111011010000101010011100101000101010101010101000101000101010100010100001000100111111111111111111111111111111111111111001000001101100111111101111111010110110000,
	240'b101100011111111111100100010110101011010011111111111111111111111111111111111111111100000001010010010100101000010111001001110000100111011101010010010100001000100111111111111111111111111111111111111111111011100001101001111101111111010110110000,
	240'b101100011111111111100100010110010111100111111001111111111111111111111111111111101000110001001100011100111111000011111111111111111110000001100011010011101000100111111111111111111111111111111111111111111110001001111001111101011111010110110000,
	240'b101100011111111111100100010111000101010111001010111111111111111111111111111101110111100001001100101000001111111111111111111111111111111110000111010010111000100111111111111111111111111111111111111111111111100110010100111100111111010110110000,
	240'b101100011111111111100100010111010100111101111111111110011111111111111111111110000111100101001100100111101111111111111111111111111111111110000101010010111000111111111111111111111111111111111111111111111111111110110110111100101111010110110000,
	240'b101100011111111111100100010111010101001101010101101111011111111111111111111111101001000001001100011011101110101011111111111111111101100001100000010011101010101011111111111111111111111111111111111111111111111111010000111101001111010110110000,
	240'b101100011111111111100100010111010101001101010010011010101110100011111111111111111100011101010100010100010111110010111101101101110110111101010000010111011101110111111111111111111111111111111111111111111111111111100100111110011111010010110000,
	240'b101100011111111111100100010111010101001101010101010100001000101011110111111111111111100110001111010011110101000001010011010100100101000001010001101001011111111011111111111111111111111111111111111111111111111111110011111111011111010010110000,
	240'b101100011111111111100100010111010101001101010101010101000101001010100010111111001111111111110001100101110101111001010100010101010110001010100111111110011111111111111111111111111111111111111111111111111111111111111010111111111111001110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010001010101101010101111110111111111111100001011111110100010101001011100011011110111111111111111111111111111111111111111111111111111111111111111111111111101111111111111001110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010100010101011010000011111000101111100111000101110101011101010111010011001111111111111111111111111111111111111111111111111111111111111111111111101111111111001111010010110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101000101001010001001110101111110100111100111111001011110010111110110111111111111111111111111111111111111111111111111111111111111111111001000111101001111010110110000,
	240'b101100011111111111100100010111010101001101010001010100010101000101010101010101010101010001010000011010101011011111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010001001111101001111010110110000,
	240'b101100011111111111100100010111010101001001111100101000000111110101010100010101010101010101010101010100100101001101110100101100011110010111111101111111111111111111111111111111111111111111111111111101001000111001101001111101111111010110110000,
	240'b101100011111111111100100010110011000101011110100111011111111010010001101010100010101010101010101010101010101010101010001010100100110010110000110101011011100011111010111110111111101110111000010011111110100111101101100111101111111010110110000,
	240'b101100011111111111100011011000001101010010111111011000111011110111011000010110000101010001010101010101010101010101010101010101010101001101010001010100000101010001011101011000010110000001010100010100010101001001101100111101111111010110110000,
	240'b101100011111111111100011011001101110010110011001010000111001100011100100010111100101001101010101010101010101010101010101010101010101010101010101010101010101010001010100010100110101001101010100010101010101001001101100111101111111010110110000,
	240'b101100011111111111100011011001101110010111100011100111111110010011000000010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100011111111111100011011001101110001011101001111010111100101001101000010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100101111111111100011011000111101110110101101011001010111011101100001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101011001111111011100110010110111010011111110100110001011110111010010110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111110001111001110101011,
	240'b100100001111100111110110011101100101010110100111110100111010011001011100010100100101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100110100110110001101111111101110100010010101,
	240'b101001111110011011111111110100000110111001011001010111100101101001011100010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010111101011100000111111111101011110100110,
	240'b111011001100001011111010111111111110111111011111110111101101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111000001111010011111111111101001100010011101010,
	240'b111111011101011111000011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111011110010011111101,
	240'b111011111111100111011110101100101011001110111101101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011000010110000110110101111001011101111,
	240'b111111111111101011100100101000001001101010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101011111001011110110100111110111111111111111111,
	240'b111111111110110010110110110101101111010111110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111001011001111110001001111100111111111,
	240'b111110111100000111100111111111111111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111111111111111111111110111001100110011111011,
	240'b110001101101011011111111111100001010100110001010100010011000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010011000011010000101100010101011010011111000111111111100110011000010,
	240'b100011111111010011111101100101100100111001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010000010100010111010110001011011000110100111010101110111111111110001110010101,
	240'b101000011111110011101011011000110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100110011111010111110100111000100110101101110010111110111110111110100010,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100100001001111001110011110111001011010101101000111101111111010110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010110101001100110101101110100011100110101101010111101111111010110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100101100101111011011100011111111111100101101101010111101111111010110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100110111011101001010101011001110010101101000001101010111101111111010110110000,
	240'b101100011111111111100100010111010101001101010011010100000101000001010000010011110101000001010010010101000101010101010101010101010101010101010101010101010101001001101011111100011000000101001001101110111100101001101010111101111111010110110000,
	240'b101100011111111111100100010111010100111101100000100010101010001010100001100101011000001101101100010110000101000001010010010101000101010101010101010101010101010001011000110010111110010010111011111101011001010101101000111101111111010110110000,
	240'b101100011111111111100100010110010111100011011000111111101111111111111111111111111111101111101110110100101010010101110010010100110101000101010101010101010101010101010010011011001100010111100000101001110101011001101011111101111111010110110000,
	240'b101100011111111111100010011100101110001111111111111111111111111111111111111111111111111111111111111111111111111111110001101110100111000101010001010101000101010101010101010100100101011001011101010100110101000101101100111101111111010110110000,
	240'b101100011111111111100000101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110100000010110000101001001010101010101010101010001010011010101010101001001101100111101111111010110110000,
	240'b101100011111110111101101111010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000100110001101010001010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100011111110011111010111101111111111111111111111111111111111111111111111111111111111111111111111111111111110011110010111100111111111011111111111111111101010001101010010100010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100011111110011111011111110011111111111111111111111111111111111111111111111111111111111111111110011101000011101101001011010111001000011011100111111111111111111011000011010000101001001010101010101010101001001101100111101111111010110110000,
	240'b101100011111110011111000111101011111111111111111111111111111111111111111111111111111111110111011010110110100111101001110010011100100111001100101110100001111111111111111110011010101110001010011010101010101001001101100111101111111010110110000,
	240'b101100011111110111110011111011101111111111111111111111111111111111111111111111111110001001011111010011100101101001111100011110010101011101001110011100011111000011111111111111111010111001010011010101010101001001101100111101111111010110110000,
	240'b101100011111111011101001111000011111111111111111111111111111111111111111111111111111000110100100011010011011110011111011111110001010110001010101010100011011110111111111111111111111100010000011010100000101001001101100111101111111010110110000,
	240'b101100011111111011100010110011011111111111111111111111111111111111111111111111111111111111111111111011001111111111111111111111111111110001110111010011001001011111111111111111111111111111011000010111000101000001101100111101111111010110110000,
	240'b101100011111111111011111101010111111111111111111111111111111111111111111111111111111111111111111111111001100111010101101101011101101011010001010010011001000101011111111111111111111111111111111100101100100110101101100111101111111010110110000,
	240'b101100011111111111100000100010011111101011111111111111111111111111111111111111111111111111101011100010100101011101010000010100000101110001011111010011111000100111111111111111111111111111111111110110100101100101101011111101111111010110110000,
	240'b101100011111111111100011011010001110001011111111111111111111111111111111111111111111011010000101010011100101000101010101010101000101000101010100010100001000100111111111111111111111111111111111111111001000001101100111111101111111010110110000,
	240'b101100011111111111100100010110101011010011111111111111111111111111111111111111111100000001010010010100101000010111001001110000100111011101010010010100001000100111111111111111111111111111111111111111111011100001101001111101111111010110110000,
	240'b101100011111111111100100010110010111100111111001111111111111111111111111111111101000110001001100011100111111000011111111111111111110000001100011010011101000100111111111111111111111111111111111111111111110001001111001111101011111010110110000,
	240'b101100011111111111100100010111000101010111001010111111111111111111111111111101110111100001001100101000001111111111111111111111111111111110000111010010111000100111111111111111111111111111111111111111111111100110010100111100111111010110110000,
	240'b101100011111111111100100010111010100111101111111111110011111111111111111111110000111100101001100100111101111111111111111111111111111111110000101010010111000111111111111111111111111111111111111111111111111111110110110111100101111010110110000,
	240'b101100011111111111100100010111010101001101010101101111011111111111111111111111101001000001001100011011101110101011111111111111111101100001100000010011101010101011111111111111111111111111111111111111111111111111010000111101001111010110110000,
	240'b101100011111111111100100010111010101001101010010011010101110100011111111111111111100011101010100010100010111110010111101101101110110111101010000010111011101110111111111111111111111111111111111111111111111111111100100111110011111010010110000,
	240'b101100011111111111100100010111010101001101010101010100001000101011110111111111111111100110001111010011110101000001010011010100100101000001010001101001011111111011111111111111111111111111111111111111111111111111110011111111011111010010110000,
	240'b101100011111111111100100010111010101001101010101010101000101001010100010111111001111111111110001100101110101111001010100010101010110001010100111111110011111111111111111111111111111111111111111111111111111111111111010111111111111001110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010001010101101010101111110111111111111100001011111110100010101001011100011011110111111111111111111111111111111111111111111111111111111111111111111111111101111111111111001110110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010100010101011010000011111000101111100111000101110101011101010111010011001111111111111111111111111111111111111111111111111111111111111111111111101111111111001111010010110000,
	240'b101100011111111111100100010111010101001101010101010101010101010101010101010101000101001010001001110101111110100111100111111001011110010111110110111111111111111111111111111111111111111111111111111111111111111111001000111101001111010110110000,
	240'b101100011111111111100100010111010101001101010001010100010101000101010101010101010101010001010000011010101011011111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010001001111101001111010110110000,
	240'b101100011111111111100100010111010101001001111100101000000111110101010100010101010101010101010101010100100101001101110100101100011110010111111101111111111111111111111111111111111111111111111111111101001000111001101001111101111111010110110000,
	240'b101100011111111111100100010110011000101011110100111011111111010010001101010100010101010101010101010101010101010101010001010100100110010110000110101011011100011111010111110111111101110111000010011111110100111101101100111101111111010110110000,
	240'b101100011111111111100011011000001101010010111111011000111011110111011000010110000101010001010101010101010101010101010101010101010101001101010001010100000101010001011101011000010110000001010100010100010101001001101100111101111111010110110000,
	240'b101100011111111111100011011001101110010110011001010000111001100011100100010111100101001101010101010101010101010101010101010101010101010101010101010101010101010001010100010100110101001101010100010101010101001001101100111101111111010110110000,
	240'b101100011111111111100011011001101110010111100011100111111110010011000000010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100011111111111100011011001101110001011101001111010111100101001101000010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101100101111111111100011011000111101110110101101011001010111011101100001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101100111101111111010110110000,
	240'b101011001111111011100110010110111010011111110100110001011110111010010110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111110001111001110101011,
	240'b100100001111100111110110011101100101010110100111110100111010011001011100010100100101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100110100110110001101111111101110100010010101,
	240'b101001111110011011111111110100000110111001011001010111100101101001011100010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010111101011100000111111111101011110100110,
	240'b111011001100001011111010111111111110111111011111110111101101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111111000001111010011111111111101001100010011101010,
	240'b111111011101011111000011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111011110010011111101,
	240'b111011111111100111011110101100101011001110111101101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011000010110000110110101111001011101111,
	240'b111111111111101011100100101000001001101010110010101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101101001011010010110100101011111001011110110100111110111111111111111111,
	240'b111111111110110010110110110101101111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111001011001111110001001111100111111111,
	240'b111110111100000111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001100110011111011,
	240'b110001101101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011000010,
	240'b100011111111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001110010101,
	240'b101000011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010100010,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101100101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110000,
	240'b101011001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110101011,
	240'b100100001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010010101,
	240'b101001111110011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011110100110,
	240'b111011001100001011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001100010011101010,
	240'b111111011101011111000011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111011110010011111101,
	240'b111011111111100111011110101100101011001110111101101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011000010110000110110101111001011101111,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule