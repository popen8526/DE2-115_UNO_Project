module yellow_eight(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111111011111110111101001100111111000100010101001101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010101000100110100011111100101111111111111101,
	240'b111111111111000110111000110110101111010011111010111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110101111010011011101101111111111001011111111,
	240'b111110011100001011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101100001011111001,
	240'b101111101101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010110111110,
	240'b100101101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010010000,
	240'b101010101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010100111,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101101011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110110011,
	240'b101001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010100011,
	240'b100101001110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110001111,
	240'b110001101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111000111,
	240'b111111011100011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101100010111111100,
	240'b111110111111001010111111110100011110111011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001110111011010010101111111111001111111011,
	240'b111011111111010111110110101011001001110010101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101001110010100010111001111111000111101111,
	240'b111111011111110111101001100111111000100010101001101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010101000100110100011111100101111111111111101,
	240'b111111111111000110111000110110101111010011111010111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110101111010111011101101111111111001011111111,
	240'b111110011100001011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101100001011111001,
	240'b101111101101010011111111111101111101000010111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011110110111100101111011100111111110111111111111101010110111110,
	240'b100101101110111111111111110010111010011010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111011100011001011101101011010010111001001111111101111010010010000,
	240'b101010101111100011111000101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101101111111001011111001111011101011000110110001111101101111100110100111,
	240'b101101011111101011110101101100011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110010001111010011000100111110001011111110101110111101001111101110110011,
	240'b101101011111101011110101101100011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111101111101011110000111110001011011010101110111101001111101110110011,
	240'b101101011111101011110101101100011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001110101011111100011100110111110011100110110101110111101001111101110110011,
	240'b101101011111101011110101101100011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100101100111110100110110101111110101110110010111100111111101110110011,
	240'b101101011111101011110101101100011010100110101001101010001010100110101001101010001010011110101000101010011010101010101010101010101010101010101010101010101010100110101111111100101100111110100110110101111110110010110010111100111111101110110011,
	240'b101101101111101011110101101100011010011110110011110011101101110011011100110110001100110111000000101100011010100110101000101010011010101010101010101010101010101010101001110101111111101011101000111110111100111010101110111101001111101110110011,
	240'b101101101111101011110101101011111011111011110001111111111111111111111111111111111111111111111101111100111101111111000011101011011010100010101010101010101010101010101001101011101101001111100100110011101010101110101111111101001111101110110011,
	240'b101101101111101011110100101111011111001111111111111111111111111111111111111111111111111111111111111111111111111111111101111010101100010010101010101010001010101010101010101010011010100010101010101010001010100110110000111101001111101110110011,
	240'b101101101111101011110100111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111101101001010100010101010101010101010101010101010101010101010100110110000111101001111101110110011,
	240'b101101101111100111111010111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001011111010101000101010101010101010101010101010101010100110110000111101001111101110110011,
	240'b101101011111100111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111101111101110111011101111101111111111111111111111011011000011101010001010101010101010101010101010100110110000111101001111101110110011,
	240'b101101011111100111111101111111101111111111111111111111111111111111111111111111111111111111111111111100001100000010101110101011101011111111101110111111111111111111111000110000101010100010101010101010101010100110110000111101001111101110110011,
	240'b101101011111100111111100111111001111111111111111111111111111111111111111111111111111111111111000101110111010011010100111101001111010011010111010111101111111111111111111111101001011100110101000101010101010100110110000111101001111101110110011,
	240'b101101011111100111111010111101011111111111111111111111111111111111111111111111111111111111011111101010001010101011000101110001101010101110100111110111001111111111111111111111111110100110101110101010011010100110110000111101001111101110110011,
	240'b101101011111100111110110111011011111111111111111111111111111111111111111111111111111111111001111101001101011100011111011111111011011100110100101110011011111111111111111111111111111111111010011101010001010100110110000111101001111101110110011,
	240'b101101011111101011110011111000011111111111111111111111111111111111111111111111111111111111010001101001101011010011110010111100111011010110100110110011111111111111111111111111111111111111111000101110001010011110110000111101001111101110110011,
	240'b101101101111101011110011110011111111111111111111111111111111111111111111111111111111111111100111101011001010100110110111101101111010100110101011111001011111111111111111111111111111111111111111110111011010100010110000111101001111101110110011,
	240'b101101101111101011110100101111101111100011111111111111111111111111111111111111111111111111101011101011111010100110100111101001111010100110101110111010011111111111111111111111111111111111111111111110011011011010101110111101001111101110110011,
	240'b101101101111101011110101101100101110011111111111111111111111111111111111111111111111100110111100101010001010100110110001101100101010101010101000101110101111100011111111111111111111111111111111111111111101001110101101111101001111101110110011,
	240'b101101101111101011110101101011101100110011111111111111111111111111111111111111111101110110101000101010011100111011110100111101011101000010101010101010001101101011111111111111111111111111111111111111111110110010110011111100111111101110110011,
	240'b101101101111101011110101101011111011001011110101111111111111111111111111111111111100011110100101101110111111101111111111111111111111110010111101101001011100010011111110111111111111111111111111111111111111101111000010111100011111101110110011,
	240'b101101011111101011110101101100011010011111010101111111111111111111111111111111101011111110100101110010111111111111111111111111111111111111001101101001011011111011111100111111111111111111111111111111111111111111010011111100011111101110110011,
	240'b101101011111101011110101101100011010100010110011111100111111111111111111111111111100001110100101110000101111111111111111111111111111111111000100101001011100001011111110111111111111111111111111111111111111111111100101111100101111101010110011,
	240'b101101011111101011110101101100011010100110101000110010101111111011111111111111111101010110100110101011011110000111111111111111111110001010101101101001101101001011111111111111111111111111111111111111111111111111110000111101001111101010110011,
	240'b101101011111101011110101101100011010100110101001101010111110000111111111111111111111001010110010101001111010111011000101110001011010111010100111101100011111000011111111111111111111111111111111111111111111111111110101111110001111101010110011,
	240'b101101011111101011110101101100011010100110101010101010001011001111101110111111111111111111011111101011011010011110100110101001101010011110101100110111011111111111111111111111111111111111111111111111111111111111111001111110111111100110110011,
	240'b101101011111101011110101101100011010100110101010101010101010100010111010111100111111111111111111111001011100000010110001101100001011111111100100111111111111111111111111111111111111111111111111111111111111111111111011111111011111100110110011,
	240'b101101101111101011110101101100011010100110101010101010101010101010101000101111001111001011111111111111111111110011110101111101011111110011111111111111111111111111111111111111111111111111111111111111111111111111111010111111001111100110110011,
	240'b101101101111101011110101101100011010100110101010101010101010101010101010101010001011011111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111101111111101010110011,
	240'b101101101111101011110101101100011010100110101010101010011010101010101010101010101010100010101111110101001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111100101111101110110011,
	240'b101101101111101011110101101100011010100010101001101011001010100110101001101010101010101010101001101010011011101111100000111110101111111111111111111111111111111111111111111111111111111111111111111111111111000010111010111100101111101110110011,
	240'b101101101111101011110101101100001010110011010101111011011101101110110001101010011010101010101010101010101010100010101010101110101101011011101101111110011111111011111111111111111111111111111111111010111011100110101110111101001111101110110011,
	240'b101101011111101011110101101011111101000111111001110111111111011011011101101010101010101010101010101010101010101010101010101010001010100010101110101110011100010111001110110100111101010011000110101100001010011110110000111101001111101110110011,
	240'b101101011111101011110101101100011110110111010101101001001100100111110110101100001010100110101010101010101010101010101010101010101010101010101001101010001010011110100111101010001010100010100111101010011010100110110000111101001111101110110011,
	240'b101101011111101011110101101100011110100111011100101010101101000111110011101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101110110011,
	240'b101101011111101011110101101011111100011011111010111011111111101111010010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101110110011,
	240'b101101011111101011110101101011111011011011110110111010011111100011000000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101110110011,
	240'b101101011111101011110101101011101011110111110111110010011111001111001010101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110000111101001111101110110011,
	240'b101001111111100011111001101100111010110111101000111110111110111110110101101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110011111101111111100110100011,
	240'b100101001110110011111111110100001010011010101111110000101011001110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011111001110111111111111001010001111,
	240'b110001101100111111111111111110101101100011000111110001101100011111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010001101100011111010111111111100111111000111,
	240'b111111011100011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101100010111111100,
	240'b111110111111001010111111110100011110111011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001110111111010010101111111111001111111011,
	240'b111011111111010111110110101011001001110010101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101001110010100010111001111111000111101111,
	240'b111111011111110111101001100111111000100010101001101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010101000100110100011111100101111111111111101,
	240'b111111111111000110111000110110101111010111111011111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110111111010111011101101111111111001011111111,
	240'b111110011100001011101000111111111111111111111110111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111101111111111111111111010101100001011111001,
	240'b101111101101010011111111111010000111001000111110001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011100100110101001110100110111111100110111111111101010110111110,
	240'b100101101110111111111101011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100101100011001000000000000001011101111111001111010110010000,
	240'b101010101111101111101001000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001101101100011101101110011000001011000010101111000111111110010100111,
	240'b101101011111110111100001000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110111101111001001110111010010011111100001011110110111111111010110011,
	240'b101101011111110111100001000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111001110111111010011111010100010011000001101110110111111111010110011,
	240'b101101011111110111100001000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111110101110110011111011000110101000001101110110111111111010110011,
	240'b101101011111110111100001000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110101110110111100000001100001101100010000011000110110101111111010110011,
	240'b101101011111110111100001000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110110000110111000000000100001111100010000011000110110101111111010110011,
	240'b101101101111110111100001000101000000000000011101011011011001011110010110100010100110100101000010000101100000000000000000000000000000000000000000000000000000000000000000100001101110111110111010111100100110110100001101110110111111111010110011,
	240'b101101101111110111100001000011100011111011010101111111111111111111111111111111111111111111111000110110101001111001001010000010100000000000000000000000000000000000000000000011000111100110101111011011010000010100010001110110111111111010110011,
	240'b101101101111110111011100001110011101101111111111111111111111111111111111111111111111111111111111111111111111111111111010110000010101000000000011000000000000000000000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101101111110011011100101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010011111000111100000000000000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101101111101011101101111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110011110100000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111100111111000111110111111111111111111111111111111111111111111111111111111111111111111111111111111010011001100110010111111001111111111111111111110010101001100000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111100111111000111111001111111111111111111111111111111111111111111111111111111111111111110100010100001000001101000011010011111111001101111111111111111111101001010001110000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111100111110101111101011111111111111111111111111111111111111111111111111111111111101001001101000000000000000000000000000000000000101111111001111111111111111111110111110010110100000000000000000000000000010010110110111111111010110011,
	240'b101101011111101011101101111000101111111111111111111111111111111111111111111111111111111110011110000000000000001001010010010101000000001100000000100101111111111111111111111111111011111000001110000000000000000000010010110110111111111010110011,
	240'b101101011111101111100011110010001111111111111111111111111111111111111111111111111111111101101111000000000010101111110011111110000010110100000000011010101111111111111111111111111111111101111100000000000000000000010010110110111111111010110011,
	240'b101101011111110011011010101001001111111111111111111111111111111111111111111111111111111101110110000000000001111111011000110111000010001000000000011100001111111111111111111111111111111111101010001010110000000000010010110110111111111010110011,
	240'b101101101111110011011001011011111111111111111111111111111111111111111111111111111111111110110111000001110000000000100101001001110000000000000110101100011111111111111111111111111111111111111111100110010000000000010010110110111111111010110011,
	240'b101101101111110111011011001111011110101111111111111111111111111111111111111111111111111111000011000011110000000000000000000000000000000000001101101111101111111111111111111111111111111111111111111011000010010100001101110110111111111010110011,
	240'b101101101111110111011111000101111011011111111111111111111111111111111111111111111110101100110101000000000000000000010110000110000000000000000000001100011110100111111111111111111111111111111111111111110111101000001011110110111111111010110011,
	240'b101101101111110111100001000011000110011111111111111111111111111111111111111111111001100000000000000000010110110111011101111000010111001100000010000000001001001011111111111111111111111111111111111111111100011000011100110110011111111010110011,
	240'b101101101111110111100001000100000001100011100000111111111111111111111111111111100101011000000000001101001111001111111111111111111111011000111000000000000101000011111101111111111111111111111111111111111111001001001000110101011111111010110011,
	240'b101101011111110111100001000100110000000010000001111111111111111111111111111110110011111000000000011001001111111111111111111111111111111101101000000000000011101111110111111111111111111111111111111111111111111101111011110100111111111010110011,
	240'b101101011111110111100001000101000000000000011011110111001111111111111111111111100100110000000000010010011111111011111111111111111111111101001101000000000100011111111011111111111111111111111111111111111111111110101111110101101111110110110011,
	240'b101101011111110111100001000101000000000000000000011000011111110011111111111111111000000000000000000010111010010111111111111111111010101000001100000000000111100111111111111111111111111111111111111111111111111111010001110111011111110110110011,
	240'b101101011111110111100001000101000000000000000000000001011010010111111111111111111101011000011000000000000000110001010000010100100000111000000000000101011101001011111111111111111111111111111111111111111111111111100010111010101111101110110011,
	240'b101101011111110111100001000101000000000000000000000000000001101111001100111111111111111110011111000010110000000000000000000000000000000000001001100110101111111111111111111111111111111111111111111111111111111111101101111100101111101010110011,
	240'b101101011111110111100001000101000000000000000000000000000000000000110010110110101111111111111111101011110100000100010100000100110100000010101100111111111111111111111111111111111111111111111111111111111111111111110010111101101111101010110011,
	240'b101101101111110111100001000101000000000000000000000000000000000000000000001101111101011111111111111111111111011011100001111000001111011011111111111111111111111111111111111111111111111111111111111111111111111111110001111101011111101010110011,
	240'b101101101111110111100001000101000000000000000000000000000000000000000000000000000010100110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111001101111110010110011,
	240'b101101101111110111100001000101000000000000000000000000000000000000000000000000000000000000010001100000001110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001110101011111110110110011,
	240'b101101101111110111100001000101000000000000000000000001110000000000000000000000000000000000000000000000000011001110100001111011111111111111111111111111111111111111111111111111111111111111111111111111111101000100101111110101111111111010110011,
	240'b101101101111110111100001000100100000100110000001110010001001010000010110000000000000000000000000000000000000000000000010001100011000010011001001111011101111110111111111111111111111111111111111110000110010111100001101110110111111111010110011,
	240'b101101011111110111100000000011100111010111101101100111101110010010011010000000100000000000000000000000000000000000000000000000000000000000001011001011100101001001101101011111010111110101010101000100010000000000010010110110111111111010110011,
	240'b101101011111110111011111000101101100011110000010000000000101110011100011000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111110111011111000101001011110010010111000010010111010011011010000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111110111100000000011100101010111110010110100001111001101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111110111100001000011110010001111100101101110111110110001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110110111111111010110011,
	240'b101101011111110111100001000011010011101011100111010111001101110101011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001110110111111111010110011,
	240'b101001111111101011101011000110110000110110111001111100101101000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111001011111101110100011,
	240'b100101001110110111111110011100100000000000010000010010010001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100111111011111001010001111,
	240'b110001101100111111111111111100011000101101011000010101000101100001011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110111000100111101111111111111100111111000111,
	240'b111111011100011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000101100010111111100,
	240'b111110111111001010111111110100011110111111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011110111111010010101111111111001111111011,
	240'b111011111111010111110110101011001001110010101110101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101001110010100010111001111111000111101111,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule