module yellow_five(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110011111100111011000100110011010000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101011011001011010111001111101001111100111111000,
	240'b111111111110110010111101110000011101010111100011111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100110111101100101110111111111000001111111111111110,
	240'b111110111011111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110000111110010111111100,
	240'b110100101101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101100001111001101,
	240'b101000101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101010100111,
	240'b101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010101111,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110111000,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010111001,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110110110,
	240'b100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010010101010,
	240'b101011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011110101011,
	240'b111001001100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001100100011100010,
	240'b111111111100101111001000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100101111101111001111111111,
	240'b111101001111101011010101101101011011100010111010101110101011101010111010101110101011101010111011101110111011101110111011101110101011101010111010101110101011101010111011101110111011101110111011101110011011010010110111111010001111010111110100,
	240'b111110011111100111011000100110011010000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101011011001011010111001111101001111100111111000,
	240'b111111111110110010111101110000011101010111100011111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100110111101100101110111111111000001111111111111110,
	240'b111110111011111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110000111110010111111100,
	240'b110100101101010011111111111111001110001011011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110101111101011111010111110110011110111111111111111101101100001111001101,
	240'b101000101111100111111101110011001010100110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110101001101101001011011010110110101101101011101111101100111111111100101110100111,
	240'b101000111111111111101110101011011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110100111100101111101111111011111111001101001111001000111111111101101010101111,
	240'b101100101111111111100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101110000001100000110111111111011001101100010111111111111111110011110111000,
	240'b101100111111111111100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011011111111001001111100001101100010111111111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110110001111101111110101111101011101000010111111111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111001111110001100110010110010101100101010101111000001111111111110100010111001,
	240'b101100111111111111100110101010101010101010101001101010001010100010101000101010001010100110101001101010101010101010101010101010101010101010101010101010101010100011000001111110001011000010100101110100011100010110111111111111111110100010111001,
	240'b101100111111111111100110101010101010100010101100101110101100001111000001101111011011001110101100101010001010100010101001101010101010101010101010101010101010100110110100111101011101110111010000111110111100010110111111111111111110100010111001,
	240'b101100111111111111100110101010001011100011100101111110101111110111111101111110111111011011101000110101011011111010101100101010001010100110101010101010101010101010101001110010001111010011111000110110011010101011000001111111111110100010111001,
	240'b101100111111111111100100101101011111000011111111111111111111111111111111111111111111111111111111111111111111110011101000110001101010110010101000101010101010101010101010101010011011001010110101101010101010011011000001111111111110100010111001,
	240'b101100111111111111100101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010110111010101010001010101010101010101010101010100110101001101010101010011111000001111111111110100010111001,
	240'b101100111111111111101111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110011001010101010101001101010101010101010101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111111000111111001111111111111111111111111111111111111111111111101111101111111011111110111111101111111011111110111111101111111100111110101101010010101011101010011010101010101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111111010111111011111111111111111111111111111111111111111111101011100001110111101101111101011111010111110101111101011111010111101110001001111011011011000101010101010100110101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111111000111111001111111111111111111111111111111111111111111100011010111010100101101001101010011010100110101001101010011110100111101011111111001111111111110100011010100010101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111110101111110101111111111111111111111111111111111111111111101011100000010111010101110101011101010111010101110111011010110101001101100011111001011111111111110111100001110101000101010101010011111000001111111111110100010111001,
	240'b101100111111111111101111111101111111111111111111111111111111111111111111111111101111101011111001111110011111100111111001111110101101110110101000101100011111001011111111111111111111000110110010101010011010011111000001111111111110100010111001,
	240'b101100111111111111101001111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001010101000101100011111001011111111111111111111111111011001101010001010011111000001111111111110100010111001,
	240'b101100111111111111100101111000011111111111111111111111111111111111111111111111111111111111111111111101101110010111011100110111011100101010101001101100011111001011111111111111111111111111111001101110101010011011000001111111111110100010111001,
	240'b101100111111111111100011110011111111111111111111111111111111111111111111111111111111111111011101101101011010100110101000101010001010100110101001101100011111001011111111111111111111111111111111110111001010011011000001111111111110100010111001,
	240'b101100111111111111100100101110101111101111111111111111111111111111111111111111111101111110101011101001111010011110101001101010011010100110101000101100011111001011111111111111111111111111111111111101111011001011000000111111111110100010111001,
	240'b101100111111111111100101101011001110101011111111111111111111111111111111111101111011011010100111101100011101001111100000111000011110000111100000111000111111101011111111111111111111111111111111111111111100101010111111111111111110100010111001,
	240'b101100111111111111100110101001111100110011111111111111111111111111111111111000101010100010101011111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111000010111111111110100010111001,
	240'b101100111111111111100110101010011011001011110011111111111111111111111111110101001010011010110111111110011111111111111111111111111111110111111000111110001111111011111111111111111111111111111111111111111111001111001011111111111110100010111001,
	240'b101100111111111111100110101010101010011111001111111111111111111111111111110101001010011010111000111110101111111111111111111111111110000110110011101111011111011011111111111111111111111111111111111111111111101111011000111111111110100010111001,
	240'b101100111111111111100110101010101010100110101111111011011111111111111111111000001010100010101100111001011111111111111111111111011100001110100100101110001111101111111111111111111111111111111111111111111111111111100101111111111110100010111001,
	240'b101100111111111111100110101010101010101010101000110000001111101111111111111101011011001110100111101101011101110111101000110010101010101010100111110100101111111111111111111111111111111111111111111111111111111111110000111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010011101010011111111111111111101101110101001101001111010100110101010101010001010011110111001111101101111111111111111111111111111111111111111111111111111111111111001111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010011010110011100000111111111111111011010110101100001010100010100111101010101011110111101111111111111111111111111111111111111111111111111111111111111111111111111100111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010101010100110101111111000111111111111111111111011111101101111010111111000111111101011111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010101010101010101000101011111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111110100010111001,
	240'b101100111111111111100110101010101010101010101010101010101010101010101010101010011010110011001111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100011111111111110100010111001,
	240'b101100111111111111100110101010101010101010101000101001111010100110101010101010101010100110101000101110101110000111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011001001111111111110100010111001,
	240'b101100111111111111100110101010101010101011000000110011011011011110101001101010101010101010101010101010001010101011000001110111111111011111111111111111111111111111111111111111111111111111111111111101001011110110111111111111111110100010111001,
	240'b101100111111111111100110101010001100111011111010111110001111001110111010101010001010101010101010101010101010101010101000101010011011011011001001110110111110100011101111111100101111000011011101101110011010010111000001111111111110100010111001,
	240'b101100111111111111100100101100011111001011010101101101011110101111011110101010001010101010101010101010101010101010101010101010101010100110100111101010011010101110101110101100011010111110101001101010001010011111000001111111111110100010111001,
	240'b101100111111111111100101101011101011111110101100101000111101101011100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011010100110101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111100101101011101100010111001001110100001111011111010011101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111100100101101111111100011111000111101101101111110101111101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111000001111111111110100010111001,
	240'b101100111111111111100100101101111111011011000100101100101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111000001111111111110100010111001,
	240'b101011101111111111100101101101111111100111100110110111111110000111000101101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111000010111111111110010110110110,
	240'b100111001111111111110011101110111101111111100111111001111110100011001000101001111010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010011011010011111111111101010010101010,
	240'b101011001111000011111111110111111011011010110001101100011011001010110001101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001100010111110111111111111100011110101011,
	240'b111001001100010111111111111111111111010111101110111011101110111011101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111100001111110111111111111010001100100011100010,
	240'b111111111100101111001000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100101111101111001111111111,
	240'b111101001111101011010101101101011011100010111010101110101011101010111010101110101011101010111011101110111011101110111011101110101011101010111010101110101011101010111011101110111011101110111011101110011011010010110111111010001111010111110100,
	240'b111110011111100111011000100110011010000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101011011001011010111001111101001111100111111000,
	240'b111111111110110010111101110000011101010111100011111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100101110111101100101110111111111000001111111111111110,
	240'b111110111011111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110000111110010111111100,
	240'b110100101101010011111111111101001010100110001011100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100010001000011110000110100011011100111111111111111101101100001111001101,
	240'b101000101111101011111010011001100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110010010000100100001001100011001111000110111111111100101010100111,
	240'b101000111111111111001100000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110110001111010011110010111101100111100101011001111111111101101110101111,
	240'b101100101111111110110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001010000110100011001000000110001101000101100111101111111111110100010111000,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101011101110100101000110000111110111111111110100110111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100010101111001011100010111000110111001000111111111111111110100110111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101111011000110011100011010000101110000100101000101111111111110100110111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100111010100001001100000000011101010101001001000000111111111110100110111001,
	240'b101100111111111110110011000000000000000000000101001100100100101001000110001110000001101000000111000000000000000000000000000000000000000000000000000000000000000000011111111000101001101001110011111100110101001000111111111111111110100110111001,
	240'b101100111111111110110011000000000010101110110000111100011111101011111000111100111110001110111100100000010011101100000111000000000000000000000000000000000000000000000000010110101101111111101010100011010000010001000101111111111110100110111001,
	240'b101100111111111110101110001000111101001111111111111111111111111111111111111111111111111111111111111111111111010110111011010101100000011100000000000000000000000000000000000000000001100000100010000000010000000001000110111111111110100110111001,
	240'b101100111111111110110001100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011001000110001000000000000000000000000000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111111001110111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000011001010000000100000000000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111111101011111101011111111111111111111111111111111111111111111111011111010011110011111100111111001111110011111100111111001111110110111100000111111000000101000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111111110001111110001111111111111111111111111111111111111111111000010100101100111010001110110011101100111011001110110011101100111010010011101110010010001011000001000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111111101011111101011111111111111111111111111111111111111111110101100000101000000000000000000000000000000000000000000000000000000000000011111101101011111111011101010000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111111100001111100001111111111111111111111111111111111111111111000000100001000110000001100010011000100110001001100110010000000000000000101011101100111111111111100110100101000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111111001110111001111111111111111111111111111111111111111111111111011111000011101110111011111110111111101111111100011001101000000000000101001101100111111111111111111101010000011010000000000000000001000110111111111110100110111001,
	240'b101100111111111110111110110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101000000000000101001101100111111111111111111111111110001101000000000000000001000110111111111110100110111001,
	240'b101100111111111110110000101001011111111111111111111111111111111111111111111111111111111111111111111000111011000010010111100110000110000000000000000101001101100111111111111111111111111111101110001100000000000001000110111111111110100110111001,
	240'b101100111111111110101010011100001111111111111111111111111111111111111111111111111111111010011001001001000000000000000000000000000000000000000000000101001101100111111111111111111111111111111111100101100000000001000101111111111110100110111001,
	240'b101100111111111110101101001100001111001011111111111111111111111111111111111111111010000000000101000000000000000000000000000000000000000000000000000101001101100111111111111111111111111111111111111001100001101001000010111111111110100110111001,
	240'b101100111111111110110001000001111011111111111111111111111111111111111111111001110010010000000000000101000111101110100011101001001010010010100011101010111111000111111111111111111111111111111111111111110110000100111110111111111110100110111001,
	240'b101100111111111110110011000000000110011011111111111111111111111111111111101010000000000000000100101000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101001000111111111111110100110111001,
	240'b101100111111111110110011000000000001011111011010111111111111111111111111011111110000000000100110111011011111111111111111111111111111100011101001111010111111110011111111111111111111111111111111111111111101110001100010111111011110100110111001,
	240'b101100111111111110110011000000000000000001110000111111111111111111111111011111010000000000101010111100001111111111111111111111111010010000100000001110001110001111111111111111111111111111111111111111111111010010001010111110101110100110111001,
	240'b101100111111111110110011000000000000000000010001110010001111111111111111101000100000000000000111101100011111111111111111111110000100101100000000001010111111001011111111111111111111111111111111111111111111111010110001111110011110100110111001,
	240'b101100111111111110110011000000000000000000000000010000111111001111111111111000000001110000000000001000001001100010111010010111110000001000000000011110101111111111111111111111111111111111111111111111111111111111010011111110111110100110111001,
	240'b101100111111111110110011000000000000000000000000000000000111110111111111111111111001001000000001000000000000000000000000000000000000000000101110111000111111111111111111111111111111111111111111111111111111111111101100111111001110100010111001,
	240'b101100111111111110110011000000000000000000000000000000000000100010100010111111111111101110000101000100110000000000000000000000100011101011001111111111111111111111111111111111111111111111111111111111111111111111110111111111011110100010111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000010000101010101111111111111111110011111001001110000110101011001110111011111111111111111111111111111111111111111111111111111111111111111111111111111001111111011110100010111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000100011001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111111001110100010111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000000000000011001110000111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101101111110101110100110111001,
	240'b101100111111111110110011000000000000000000000000000000000000000000000000000000000000000000000000001100101010011011110110111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101011101111111011110100110111001,
	240'b101100111111111110110011000000000000000101000010011010000010011100000000000000000000000000000000000000000000001001000110100111111110011011111111111111111111111111111111111111111111111111111111110111110011101001000000111111111110100110111001,
	240'b101100111111111110110011000000000110110111110000111010001101110000110001000000000000000000000000000000000000000000000000000000000010010101011110100100101011101011010000110101111101001010011011001011100000000001000110111111111110100110111001,
	240'b101100111111111110110000000101001101100110000001001001101100001110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001011000101000000111000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111110110001000010110011111100000111000000001001000010110111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111110110001000011010101000101011111011100111110011101111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111110101110001001101110101111101010111000111001111100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101100111111111110101110001010001110001001001111000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110111111111110100110111001,
	240'b101011101111111110110001001010011110110110110110100111111010011001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000111111111110011010110110,
	240'b100111001111111111011001001100101001111010110110101101111011100101011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100111111111101010010101010,
	240'b101011001111000011111111100111100010010000010110000101110001011100010100000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000101000101000011100111111111111100011110101011,
	240'b111001001100010111111111111111111110000011001100110011011100110111001110110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001110110100111111011111111111111010001100100011100010,
	240'b111111111100101111001000111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100101111101111001111111111,
	240'b111101001111101011010101101101011011100010111010101110101011101010111010101110101011101010111011101110111011101110111011101110101011101010111010101110101011101010111011101110111011101110111011101110011011010010110111111010001111010111110100,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule