module yellow_nine(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111110101111110011101100101001001000111010101010101011011010110110101101101011011010110110101100101011001010110010101100101011001010110110101101101011011010110110101101101011001010110010101101101010101000111010101010111100101111110011111010,
	240'b111111111111101111000010110001101101111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111011001000110011001111110111111111,
	240'b111111111100110011010110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011100111111111110,
	240'b110010101100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100011001100,
	240'b100111011110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110010110,
	240'b101011001111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010101001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111010,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101110001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111001,
	240'b101011001111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110101001,
	240'b100110111110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010010100,
	240'b110010111100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111001100,
	240'b111111111100110111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001101000011111110,
	240'b111110101111011111000111110010011110010011100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110001111000110110010001111011111111010,
	240'b111011111111001011110110101011111010000010110101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011001111110101000111010011111000011101111,
	240'b111110101111110011101100101001001000111010101010101011011010110110101101101011011010110110101100101011001010110010101100101011001010110110101101101011011010110110101101101011001010110010101101101010101000111010101010111100101111110011111010,
	240'b111111111111101111000010110001101101111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111011001000110011001111110111111111,
	240'b111111111100110011010110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011100111111111110,
	240'b110010101100100111111111111111011110000011001110110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110011001011110011011110000111111101111111111100100011001100,
	240'b100111011110010111111111110101111010100110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001101011001110111101101011101010100011011001111111111110100010010110,
	240'b101011001111010111111100101110001010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110001001111010111111011111011011011010010111000111111001111000010101001,
	240'b101110001111110011110111101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101110111011101110000010111110111011111101101010110100111110011111001010111001,
	240'b101110001111110011110111101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111101011100000010100000110101101110100010110110111110011111001010111001,
	240'b101110001111110011110111101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110001110001111000100111100101101100010110100111110011111001010111001,
	240'b101110001111110011110111101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111101011111100111111010111001111011001010110100111110011111001010111001,
	240'b101110001111110011110111101101001010100110101001101010001010100010101000101010001010100010101000101010011010101010101010101010101010101010101010101010101010100110110011111101001100110110110110101110001010101010110101111110011111001010111001,
	240'b101110011111110011110111101101001010011110101110110000111101000111010001110011011100001010110111101011001010100010101000101010101010101010101010101010101010101010101010111000101111001111011011111100111011111110110011111110011111001010111010,
	240'b101110011111110011110111101100101011011011101000111111101111111111111111111111111111111111111000111010101101010010111010101010101010100010101010101010101010101010101001101101001110000011101101110101001010110010110101111110011111001010111010,
	240'b101110011111110011110110101110101110101111111111111111111111111111111111111111111111111111111111111111111111111111111001111000001011101110101001101010011010101010101010101010011010101010101101101010011010100010110101111110011111001010111010,
	240'b101110011111110011110101110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111010100101011101010100010101010101010101010101010101001101010101010100110110101111110011111001010111010,
	240'b101110011111101111111001111101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011011010101000101010101010101010101010101010101010100110110101111110011111001010111010,
	240'b101110001111101111111011111111011111111111111111111111111111111111111111111111111111111111111111111111111111110011110011111100111111110111111111111111111111000010111010101010001010101010101010101010101010100110110101111110011111001010111010,
	240'b101110001111101111111011111111001111111111111111111111111111111111111111111111111111111111111111111001001011111110110010101100101011111111100110111111111111111111110010101110011010100010101010101010101010100110110101111110011111001010111001,
	240'b101110001111101111111011111111001111111111111111111111111111111111111111111111111111111111011101101011001010011110100110101001101010011110101100110111101111111111111111111011011011001010101001101010101010100110110101111110011111001010111001,
	240'b101110001111101111111001111101111111111111111111111111111111111111111111111111111111000110110001101001111010111111000110110001011010111110100111101100101111001011111111111111111110000010101011101010011010100110110101111110011111001010111001,
	240'b101110001111101111110111111011011111111111111111111111111111111111111111111111111101010010100110101011011110001111111111111111111110001010101101101001111101011011111111111111111111111011001010101010001010100110110101111110011111001010111001,
	240'b101110001111110011110101111000001111111111111111111111111111111111111111111111111100001110100101110001001111111111111111111111111111111111000001101001011100010111111111111111111111111111110010101100101010011110110101111110011111001010111001,
	240'b101110011111110011110101110100001111111011111111111111111111111111111111111111101011110110100101110011001111111111111111111111111111111111001001101001011100001011111110111111111111111111111111110101001010011010110101111110011111001010111010,
	240'b101110011111110011110110110000001111011111111111111111111111111111111111111111101011110110100110101110101111101011111111111111111111100110111001101001011100101011111111111111111111111111111111111100111011000010110100111110011111001010111010,
	240'b101110011111110011110111101101001110010111111111111111111111111111111111111111101011110110101000101010011100101111110000111100001100101010101001101010011110000111111111111111111111111111111111111111111100100110110011111110011111001010111010,
	240'b101110011111110011110111101100011100101011111111111111111111111111111111111111101011110110101000101010011010100110110000101100001010100010100111110000001111101111111111111111111111111111111111111111111110010010110110111110011111001010111010,
	240'b101110011111110011110111101100101011000111110100111111111111111111111111111111101011110110101000101011001010100110100111101001111010100010111101111100101111111111111111111111111111111111111111111111111111011011000001111110001111001010111010,
	240'b101110001111110011110111101101001010011111010100111111111111111111111111111111101011110110100110110001111101110111001001110010101101110111111001111111111111111111111111111111111111111111111111111111111111111011010000111101111111001010111001,
	240'b101110001111110011110111101101001010011110110010111100101111111111111111111111111100001110100101110001001111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111100001111101111111001010111001,
	240'b101110001111110011110111101101001010100110101000110010011111111011111111111111111101010110100110101011101110001111111111111111111101111110111101111000011111110011111111111111111111111111111111111111111111111111101110111110001111001010111001,
	240'b101110001111110011110111101101001010100110101001101010111110000011111111111111111111000110110001101001111010111111000111110001011010111010100110101101001111010111111111111111111111111111111111111111111111111111110100111110101111001010111001,
	240'b101110001111110011110111101101001010100110101010101010011011001011101101111111111111111111011110101011001010011010100110101001101010011110101101110111101111111111111111111111111111111111111111111111111111111111110111111111001111000110111001,
	240'b101110001111110011110111101101001010100110101010101010101010100010111010111100111111111111111111111001101100001110110011101100111100000111100101111111111111111111111111111111111111111111111111111111111111111111111001111111011111000110111010,
	240'b101110011111110011110111101101001010100110101010101010101010101010101000101111001111000111111111111100101101011111010000110100001101011111110011111111111111111111111111111111111111111111111111111111111111111111111001111111011111000110111010,
	240'b101110011111110011110111101101001010100110101010101010101010101010101010101010001011011111101010111010001100010011000101110001011100010011101000111111111111111111111111111111111111111111111111111111111111111111110010111110011111001010111010,
	240'b101110011111110011110111101101001010100110101010101010011010101010101010101010101010100010101111110101001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010111101111111001010111010,
	240'b101110011111110011110111101101001010100010101001101011011010101010101001101010101010101010101001101010011011101011011111111110101111111111111111111111111111111111111111111111111111111111111111111111111110100110111011111110001111001010111010,
	240'b101110011111110011110111101100111010110111010101111011101101111010110011101010011010101010101010101010101010100010101010101110011101010111101100111110001111111011111111111111111111111111111101111001101011010010110100111110011111001010111010,
	240'b101110001111110011110111101100011100000111110011110110111111001111100000101010101010101010101010101010101010101010101010101010001010100010101101101110001100001111001100110100011101000111000010101011011010011110110101111110011111001010111001,
	240'b101110001111110011110111101100111010101010111001101110001100111011110101101100011010100110101010101010101010101010101010101010101010101010101001101010001010011110100111101010001010100010101000101010011010100110110101111110011111001010111001,
	240'b101110001111110011110111101100101011001111101000111110011111011111110111101100101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110011111001010111001,
	240'b101110001111110011110111101100101101101011110000110001001110010011111000101100101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110011111001010111001,
	240'b101110001111110011110111101101001110101111010100101000001100000111110111101100101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110011111001010111001,
	240'b101110001111110011110111101100101101110111101110101111111110001011101101101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110011111001010111001,
	240'b101011001111010011111100101101101011010111101110111110101111010111000010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111001111000010101001,
	240'b100110111110010011111111110101111010100010101110101111011011001110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111010100111011001111111111110011010010100,
	240'b110010111100100111111111111111011110000011001110110011011100111011001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111110000111111110111111111100011111001100,
	240'b111111111100110111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001101000011111110,
	240'b111110101111011111000111110010011110010011100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110010011000110110010001111011111111010,
	240'b111011111111001011110110101011111010000010110101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011001111110101000111010011111000011101111,
	240'b111110101111110011101100101001001000111010101010101011011010110110101101101011011010110110101100101011001010110010101100101011001010110110101101101011011010110110101101101011001010110010101101101010101000111010101010111100101111110011111010,
	240'b111111111111101111000010110001101101111111101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111011001000110011001111110111111111,
	240'b111111111100110011010110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011100111111111110,
	240'b110010101100100111111111111110011010001001101100011010010110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110011001100010011010011010010011111010111111111100100011001100,
	240'b100111011110010111111111100010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111010000011000000000010001101111111111110100010010110,
	240'b101011001111011011110011001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011011110000111110010110010000010000000101011111101001111001010101001,
	240'b101110001111111011100110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110011001010000100111110110011111001000100011100111010011111010010111001,
	240'b101110001111111011100110000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111000100100001100000000100001001011101000100011111010011111010010111001,
	240'b101110001111111011100110000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111010101010101001010000110101111000101000011101111010101111010010111001,
	240'b101110001111111011100110000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111000111110110111110001101101110001100100011110111010101111010010111001,
	240'b101110001111111011100110000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110111110110100100100101001010100000010100100001111010101111010010111001,
	240'b101110011111111011100110000111010000000000001100010011000111010101110110011010010100100100101000000001110000000000000000000000000000000000000000000000000000000000000011101010001101101010010100110110100011111100011011111010101111010010111010,
	240'b101110011111111011100110000110000010010110111001111111011111111111111111111111111111111111101010110000010111111000101111000000000000000000000000000000000000000000000000000111011010000111001010011111100000101000100000111010101111010010111010,
	240'b101110011111111011100011001100011100001111111111111111111111111111111111111111111111111111111111111111111111111111101101101000110011010000000000000000000000000000000000000000000000000000001000000000000000000000100010111010101111010010111010,
	240'b101110011111111011100000100100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001111110000011100000000000000000000000000000000000000000000000000000000000100010111010101111010010111010,
	240'b101110011111110011101011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010010011000000000000000000000000000000000000000000000000000100010111010101111010010111010,
	240'b101110001111110011110011111110001111111111111111111111111111111111111111111111111111111111111111111111111111011111011100110111001111100011111111111111111101000100110010000000000000000000000000000000000000000000100010111010101111010010111010,
	240'b101110001111110011110011111110001111111111111111111111111111111111111111111111111111111111111111101011110100000000011001000110010100001010110010111111111111111111010111001011100000000000000000000000000000000000100010111010101111010010111001,
	240'b101110001111110011110010111101101111111111111111111111111111111111111111111111111111111110011000000010010000000000000000000000000000000000001011100111011111111111111111110010100001101000000000000000000000000000100010111010101111010010111001,
	240'b101110001111110011101110111001101111111111111111111111111111111111111111111111111101010100010110000000000001000001010100010100100000111100000000000110001101100011111111111111111010001000000101000000000000000000100010111010101111010010111001,
	240'b101110001111110111100110110010011111111111111111111111111111111111111111111111111000000000000000000011001010110011111111111111111010011100001011000000001000010011111111111111111111110001011111000000000000000000100010111010101111010010111001,
	240'b101110001111111011011111101001001111111111111111111111111111111111111111111111110100110000000000010011011111111111111111111111111111111101000110000000000101000111111110111111111111111111011001000110010000000000100010111010101111010010111001,
	240'b101110011111111011011111011100011111110011111111111111111111111111111111111111010011101100000000011001011111111111111111111111111111111101011101000000000100100011111100111111111111111111111111011111010000000000100010111010101111010010111010,
	240'b101110011111111011100010010000011110011111111111111111111111111111111111111111010011101000000000001100011111000011111111111111111110111000101100000000000110000011111111111111111111111111111111110111000001001100011110111010101111010010111010,
	240'b101110011111111011100101000111101011000111111111111111111111111111111111111111010011101000000000000000010110001111010011110100100101111100000000000000001010011011111111111111111111111111111111111111110101111000011010111010101111010010111010,
	240'b101110011111111011100110000101010110000111111111111111111111111111111111111111010011101000000000000000000000000000010011000100110000000000000000010000101111001011111111111111111111111111111111111111111010111000100011111010011111010010111010,
	240'b101110011111111011100110000110010001010011011101111111111111111111111111111111010011101000000000000001110000000000000000000000000000000000111010110101111111111111111111111111111111111111111111111111111110010101000100111001101111010010111010,
	240'b101110001111111011100110000111010000000001111101111111111111111111111111111111010011101100000000010101101001100101011101011000001001100111101101111111111111111111111111111111111111111111111111111111111111110001110011111000111111010010111001,
	240'b101110001111111011100110000111010000000000011001110110101111111111111111111111110100110000000000010011101111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111110100101111000111111010010111001,
	240'b101110001111111011100110000111010000000000000000010111101111101111111111111111111000000000000000000011011010110011111111111111111001111100111011101001001111011111111111111111111111111111111111111111111111111111001011111001011111010010111001,
	240'b101110001111111011100110000111010000000000000000000001001010001111111111111111111101011000010111000000000000111101010110010100110000101100000000000111011110001011111111111111111111111111111111111111111111111111011110111011011111001110111001,
	240'b101110001111111011100110000111010000000000000000000000000001101011001010111111111111111110011100000010100000000000000000000000000000000000001010100111011111111111111111111111111111111111111111111111111111111111101000111101001111001010111001,
	240'b101110001111111011100110000111010000000000000000000000000000000000110000110110101111111111111111101100100100101100011011000110100100011110110010111111111111111111111111111111111111111111111111111111111111111111101101111101111111001010111010,
	240'b101110011111111011100110000111010000000000000000000000000000000000000000001101101101011011111111110110001000011101110010011100011000011011011010111111111111111111111111111111111111111111111111111111111111111111101101111101101111001010111010,
	240'b101110011111111011100110000111010000000000000000000000000000000000000000000000000010100011000001101110100100111101010010010100100100110110111010111111111111111111111111111111111111111111111111111111111111111111011001111010111111001110111010,
	240'b101110011111111011100110000111010000000000000000000000000000000000000000000000000000000000010000011111101110101111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111110010000111000111111010010111010,
	240'b101110011111111011100110000111010000000000000000000010010000000000000000000000000000000000000000000000000011001110100001111011111111111111111111111111111111111111111111111111111111111111111111111111111011110000110010111010001111010010111010,
	240'b101110011111111011100110000110110000101110000001110010111001110000011010000000000000000000000000000000000000000000000001001011101000000111000101111010111111110011111111111111111111111111111010101100110010000000011101111010101111010010111010,
	240'b101110001111111011100110000101110100010111011011100100111101101110100001000000110000000000000000000000000000000000000000000000000000000000001001001010100100110001100110011101100111010001001001000010010000000000100010111010101111010010111001,
	240'b101110001111111011100110000111000000010100101100001011010110110011100010000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111010101111010010111001,
	240'b101110001111111011100110000110010001110010111010111010111110100011100111000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111010101111010010111001,
	240'b101110001111111011100110000110001001000111010011010100101010111011101100000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111010101111010010111001,
	240'b101110001111111011100101000111011100001101111101000000000100010111101000000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111010101111010010111001,
	240'b101110001111111011100110000101111001100011001011010000101010011111001000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111010101111010010111001,
	240'b101011001111011011110011001001010010001011001100111100001110000101000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111101001111001010101001,
	240'b100110111110010111111111100010000000000000001101001110010001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001101111111111110011010010100,
	240'b110010111100100011111111111110011010001001101100011010000110101101101110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110011011111010010111111010111111111100011111001100,
	240'b111111111100110111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001101000011111110,
	240'b111110101111011111000111110010011110010011100111111010001110011111100111111001111110011111100111111010001110100011101000111010001110011111100111111001111110011111100111111010001110100011101000111001111110010011000110110010001111011111111010,
	240'b111011111111001011110110101011111010000010110101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011001111110101000111010011111000011101111,
};
assign data = picture[addr];
endmodule