module red_six(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111011111111011111101100110000011011000110110010101100111011001010110010101100101011001010110011101100111011001110110011101100111011001010110010101100101011001010110011101100111011001110110011101100111011000011000000111001101111000111101111,
	240'b111100011110011010111111110111101111100011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111011111011010101110001110000111110010,
	240'b111001111011110011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011101011101001,
	240'b101100111101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011110110100,
	240'b100100001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001101,
	240'b101010001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110100010,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110000,
	240'b101101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110001,
	240'b101011001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010100110,
	240'b100100011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110001101,
	240'b101010101110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111010101010,
	240'b111000011011110111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011011110011100011,
	240'b111100101101101111000001111011101111111111111110111111011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111101111111101111111111101011101110101101100011110010,
	240'b111110011111101011011110100111011001101010101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001100010100101111001101111110011111001,
	240'b111011111111011111101100110000101011000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011000111000000111001101111000111101111,
	240'b111100011110011010111111110111101111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111100011011010101110001110000111110010,
	240'b111001111011110011110000111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111011001011101011101001,
	240'b101100111101110011111111111010001001101001111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111101001111000011110101001111011101101111111111101011110110100,
	240'b100100001111110011111001100001100100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010111011110011000011100110100101110010000111111001111011010001101,
	240'b101010001111111111100001010111000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100100001111010111101111111100011000010001011101111010111111111010100010,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011111101001101001101000110000111101001001011101111001011111111110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110011001110010111100110010101110001001100011111001011111111110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101010101111011011010110111110101110001001100011111001011111111110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001111010000101001111101011101110011001100011111001011111111110110000,
	240'b101101101111111111011011010110010101010001010011010100000101001001010010010100000101000001010001010100110101010101010101010101010101010101010101010101010101001101011111111010011001101001001011101010001101111001100001111001011111111110110000,
	240'b101101101111111111011011010110010101000001101000100110101011000010101111101001111001001101111010011000000101001001010001010101000101010101010101010101010101010101010011101101001111001011000111111101011010011001011001111001101111111110110000,
	240'b101101101111111111011011010101011000011111100100111111111111111111111111111111111111111111110111111000011011100010000000010101110101000101010100010101010101010101010011011000001010111011010010101001110101101101011011111001101111111110110000,
	240'b101101101111111111010111011110101110111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010101000000001010011010100100101010101010101010100110101001101010111010100100101001101011100111001101111111110110000,
	240'b101101101111111111011010110001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110100011000110101000101010101010101010101010101010100010101010101010001011100111001101111111110110000,
	240'b101101101111111111101100111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111010101010000010101010101010101010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111111001111110011111111111111111111111111111111111111111111111111111111111111111111111111111011111100110111010001111100111111111111111111110100001111110010100000101010101010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111111010111110101111111111111111111111111111111111111111111111111111111111111110110000100111101101011111011000000111111111001011111111111111111111101011011110100101000001010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111110110111101101111111111111111111111111111111111111111111111111111111010110000010101100100111101001110010011100100111001011010101111001111111111111111111000100110101101010001010101010101010001011100111001101111111110110000,
	240'b101101101111111111101111111011111111111111111111111111111111111111111111111111111110000101011101010011010101111010001001100010010101110101001111011000111110001111111111111111111100100101011001010101000101010001011100111001101111111110110000,
	240'b101101101111111111100011111001001111111111111111111111111111111111111111111111111111011010110100011101001100010011111111111111111100000101011010010011101010100111111111111111111111111110011110010100010101001101011100111001101111111110110000,
	240'b101101101111111111011011110100001111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111110000101010011001000011111111101111111111111111111101100011011000101000001011100111001101111111110110000,
	240'b101101101111111111010110101011011111111111111111111111111111111111111111111111111111111111111111111101011100000010011010100110111100010110010000010011010111110011111010111111111111111111111111101101000101000001011100111001101111111110110000,
	240'b101101101111111111010110100010011111110011111111111111111111111111111111111111111111111111100010011111000101001101001110010011110101011001011100010100010111110011111010111111111111111111111111111011110110101001011001111001101111111110110000,
	240'b101101101111111111011001011001101110010111111111111111111111111111111111111111111111001101111100010011100101000101011100010110110101000101010100010100010111110011111010111111111111111111111111111111111010000101010111111001101111111110110000,
	240'b101101101111111111011011010101101011011011111111111111111111111111111111111111111011100101010001010100111001000111011001110101101000101001010011010100010111110011111010111111111111111111111111111111111101011001100001111001011111111110110000,
	240'b101101101111111111011011010101000111101011111001111111111111111111111111111111011000100101001100011101111111010111111111111111111110111101101111010011100111110011111010111111111111111111111111111111111111010101111110111000101111111110110000,
	240'b101101101111111111011011010110000101010111001000111111111111111111111111111101110111011101001100100111111111111111111111111111111111111110010100010011000111110011111010111111111111111111111111111111111111111110100001111000011111111110110000,
	240'b101101101111111111011011010110010100111101111100111110001111111111111111111110010111101101001100100101011111111111111111111111111111111110001011010011001000010011111101111111111111111111111111111111111111111111000100111000101111111110110000,
	240'b101101101111111111011011010110010101001101010011101101101111111111111111111111111001011001001101011001011101110011111111111111111101010101100000010011011010000111111111111111111111111111111111111111111111111111011100111010011111111110110000,
	240'b101101101111111111011011010110010101010001010010011001001110000011111111111111111101000001011000010100000110110010100111101001000110100001010000010111001101100111111111111111111111111111111111111111111111111111101100111100111111111010110000,
	240'b101101101111111111011011010110010101010001010101010100010111111011110001111111111111110110100001010100100100111101010000010100000100111101010011101010101111111011111111111111111111111111111111111111111111111111110110111110101111111010110000,
	240'b101101101111111111011011010110010101010001010101010101010101000110010010111101111111111111111010101011110110110001011011010110110110111110110110111111001111111111111111111111111111111111111111111111111111111111111011111111011111110110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010001010010100101111111011011111111111011011011111110100101101001101100000111110001111111111111111111111111111111111111111111111111111111111111111111111101111111101111110110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010100010100101000101111101111110001000111010101111001011110010111010111000111111111111111111111111111111111111111111111111111111111111111111111110000111101011111111010110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101000101000101110111110010101111010011110110111100111111001011111010111111111111111111111111111111111111111111111111111111111111111111001001111001011111111110110000,
	240'b101101101111111111011011010110010101001101010001010100100101000101010100010101010101010101010001010111011001110011100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010000010111000101111111110110000,
	240'b101101101111111111011011010110000101011110010011101101111000111101010110010101000101010101010101010100110101000001100100100110011101001011110100111111111111111111111111111111111111111111111111111100001001000001011001111001101111111110110000,
	240'b101101101111111111011011010101011001111111111000111000101111011110011000010100010101010101010101010101010101010101010011010100000101100101110001100101001010111011000010110011001100110110110001011101010101000001011100111001101111111110110000,
	240'b101101101111111111011001011000011110000010101011010101001011001111011100010110010101010001010101010101010101010101010101010101010101010001010010010100000101000001010101010110000101100001010010010100010101010001011100111001101111111110110000,
	240'b101101101111111111011001011001101110101110010111010001111010001011100010010111000101001101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111011001011001101110101111101100101110101111000010110000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111011001011001101110100011010111110110101011000001011110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111001101111111110110000,
	240'b101101111111111111011001011000001110000010101101011000101000011001101011010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111001101111111110110001,
	240'b101011001111111111011111010110001001111111110110110111101111010110001111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111010011111111010100110,
	240'b100100011111110111110101011110010101000010010000101101101000101001010101010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100110110000010111110011111100010001101,
	240'b101010101110010011111111110110010111111101100110011001110110011101101010011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010101000010011100000111111111101111010101010,
	240'b111000011011110111111000111111111111100111110000111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111101011111111111101011011110011100011,
	240'b111100101101101111000001111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011101110101101100011110010,
	240'b111110011111101011011110100111011001101010101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001100010100101111001101111110011111001,
	240'b111011111111011111101100110000011011000110110010101100111011001010110010101100101011001010110011101100111011001110110011101100111011001010110010101100101011001010110011101100111011001110110011101100111011000011000000111001101111000111101111,
	240'b111100011110011010111111110111101111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111100011011010101110001110000111110010,
	240'b111001111011110011110000111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111011001011101011101001,
	240'b101100111101110011111111111010001001101001111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111101001111000011110101001111011101101111111111101011110110100,
	240'b100100001111110011111001100001100100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010111011110011000011100110100101110010000111111001111011010001101,
	240'b101010001111111111100001010111000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100100001111010111101111111100011000010001011101111010111111111010100010,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011111101001101001101000110000111101001001011101111001011111111110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110011001110010111100110010101110001001100011111001011111111110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101010101111011011010110111110101110001001100011111001011111111110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001111010000101001111101011101110011001100011111001011111111110110000,
	240'b101101101111111111011011010110010101010001010011010100000101001001010010010100000101000001010001010100110101010101010101010101010101010101010101010101010101001101011111111010011001101001001011101010001101111001100001111001011111111110110000,
	240'b101101101111111111011011010110010101000001101000100110101011000010101111101001111001001101111010011000000101001001010001010101000101010101010101010101010101010101010011101101001111001011000111111101011010011001011001111001101111111110110000,
	240'b101101101111111111011011010101011000011111100100111111111111111111111111111111111111111111110111111000011011100010000000010101110101000101010100010101010101010101010011011000001010111011010010101001110101101101011011111001101111111110110000,
	240'b101101101111111111010111011110101110111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010101000000001010011010100100101010101010101010100110101001101010111010100100101001101011100111001101111111110110000,
	240'b101101101111111111011010110001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110100011000110101000101010101010101010101010101010100010101010101010001011100111001101111111110110000,
	240'b101101101111111111101100111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111010101010000010101010101010101010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111111001111110011111111111111111111111111111111111111111111111111111111111111111111111111111011111100110111010001111100111111111111111111110100001111110010100000101010101010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111111010111110101111111111111111111111111111111111111111111111111111111111111110110000100111101101011111011000000111111111001011111111111111111111101011011110100101000001010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111110110111101101111111111111111111111111111111111111111111111111111111010110000010101100100111101001110010011100100111001011010101111001111111111111111111000100110101101010001010101010101010001011100111001101111111110110000,
	240'b101101101111111111101111111011111111111111111111111111111111111111111111111111111110000101011101010011010101111010001001100010010101110101001111011000111110001111111111111111111100100101011001010101000101010001011100111001101111111110110000,
	240'b101101101111111111100011111001001111111111111111111111111111111111111111111111111111011010110100011101001100010011111111111111111100000101011010010011101010100111111111111111111111111110011110010100010101001101011100111001101111111110110000,
	240'b101101101111111111011011110100001111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111110000101010011001000011111111101111111111111111111101100011011000101000001011100111001101111111110110000,
	240'b101101101111111111010110101011011111111111111111111111111111111111111111111111111111111111111111111101011100000010011010100110111100010110010000010011010111110011111010111111111111111111111111101101000101000001011100111001101111111110110000,
	240'b101101101111111111010110100010011111110011111111111111111111111111111111111111111111111111100010011111000101001101001110010011110101011001011100010100010111110011111010111111111111111111111111111011110110101001011001111001101111111110110000,
	240'b101101101111111111011001011001101110010111111111111111111111111111111111111111111111001101111100010011100101000101011100010110110101000101010100010100010111110011111010111111111111111111111111111111111010000101010111111001101111111110110000,
	240'b101101101111111111011011010101101011011011111111111111111111111111111111111111111011100101010001010100111001000111011001110101101000101001010011010100010111110011111010111111111111111111111111111111111101011001100001111001011111111110110000,
	240'b101101101111111111011011010101000111101011111001111111111111111111111111111111011000100101001100011101111111010111111111111111111110111101101111010011100111110011111010111111111111111111111111111111111111010101111110111000101111111110110000,
	240'b101101101111111111011011010110000101010111001000111111111111111111111111111101110111011101001100100111111111111111111111111111111111111110010100010011000111110011111010111111111111111111111111111111111111111110100001111000011111111110110000,
	240'b101101101111111111011011010110010100111101111100111110001111111111111111111110010111101101001100100101011111111111111111111111111111111110001011010011001000010011111101111111111111111111111111111111111111111111000100111000101111111110110000,
	240'b101101101111111111011011010110010101001101010011101101101111111111111111111111111001011001001101011001011101110011111111111111111101010101100000010011011010000111111111111111111111111111111111111111111111111111011100111010011111111110110000,
	240'b101101101111111111011011010110010101010001010010011001001110000011111111111111111101000001011000010100000110110010100111101001000110100001010000010111001101100111111111111111111111111111111111111111111111111111101100111100111111111010110000,
	240'b101101101111111111011011010110010101010001010101010100010111111011110001111111111111110110100001010100100100111101010000010100000100111101010011101010101111111011111111111111111111111111111111111111111111111111110110111110101111111010110000,
	240'b101101101111111111011011010110010101010001010101010101010101000110010010111101111111111111111010101011110110110001011011010110110110111110110110111111001111111111111111111111111111111111111111111111111111111111111011111111011111110110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010001010010100101111111011011111111111011011011111110100101101001101100000111110001111111111111111111111111111111111111111111111111111111111111111111111101111111101111110110110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010100010100101000101111101111110001000111010101111001011110010111010111000111111111111111111111111111111111111111111111111111111111111111111111110000111101011111111010110000,
	240'b101101101111111111011011010110010101010001010101010101010101010101010101010101000101000101110111110010101111010011110110111100111111001011111010111111111111111111111111111111111111111111111111111111111111111111001001111001011111111110110000,
	240'b101101101111111111011011010110010101001101010001010100100101000101010100010101010101010101010001010111011001110011100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010000010111000101111111110110000,
	240'b101101101111111111011011010110000101011110010011101101111000111101010110010101000101010101010101010100110101000001100100100110011101001011110100111111111111111111111111111111111111111111111111111100001001000001011001111001101111111110110000,
	240'b101101101111111111011011010101011001111111111000111000101111011110011000010100010101010101010101010101010101010101010011010100000101100101110001100101001010111011000010110011001100110110110001011101010101000001011100111001101111111110110000,
	240'b101101101111111111011001011000011110000010101011010101001011001111011100010110010101010001010101010101010101010101010101010101010101010001010010010100000101000001010101010110000101100001010010010100010101010001011100111001101111111110110000,
	240'b101101101111111111011001011001101110101110010111010001111010001011100010010111000101001101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111011001011001101110101111101100101110101111000010110000010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111001101111111110110000,
	240'b101101101111111111011001011001101110100011010111110110101011000001011110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111001101111111110110000,
	240'b101101111111111111011001011000001110000010101101011000101000011001101011010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111001101111111110110001,
	240'b101011001111111111011111010110001001111111110110110111101111010110001111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111010011111111010100110,
	240'b100100011111110111110101011110010101000010010000101101101000101001010101010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100110110000010111110011111100010001101,
	240'b101010101110010011111111110110010111111101100110011001110110011101101010011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010101000010011100000111111111101111010101010,
	240'b111000011011110111111000111111111111100111110000111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111101011111111111101011011110011100011,
	240'b111100101101101111000001111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011101110101101100011110010,
	240'b111110011111101011011110100111011001101010101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001100010100101111001101111110011111001,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule