module yellow_one(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110011111011011100011100110011001001010101011101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010111001000010100100111011111111110011111001,
	240'b111111011110100010111100110010101110000011101100111011101110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101110111011001101111011001001110010101111101111111100,
	240'b111110101011110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011100101011111101,
	240'b110010111101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011001011,
	240'b101001001111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110011100,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010101011,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110010,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110101111,
	240'b101001001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011101,
	240'b101101111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010110100,
	240'b111100011011100111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100000111110100,
	240'b111111011101110010111011111001111111110111111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011100001101111001110110111111101,
	240'b111101001111111111101010101011001010000110101001101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101011101010111010101110101011101010011001111110101010111001011111001111110100,
	240'b111110011111011011100011100110011001001010101011101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010111001000010100100111011111111110011111001,
	240'b111111011110100010111100110010101110000011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111011001001110010101111101111111100,
	240'b111110101011110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011100101011111101,
	240'b110010111101000111111111111110111101110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001110110011011110000011111101111111111100110011001011,
	240'b101001001111010011111110110011101010100010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110110101101110001010100011010101111111111110110110011100,
	240'b101011101111111111110100101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011011100111110111100010010110101111110011111100110101011,
	240'b101101001111111111101101101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011011101111101111110010010110101111101001111100110110010,
	240'b101101001111111111101101101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011011110111000001011110010110101111101001111101010110010,
	240'b101101001111111111101101101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011011110110111111010011110110010111101001111101010110010,
	240'b101101001111111111101101101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011011110110111111010100010110010111101001111101010110010,
	240'b101101001111111111101101101011101010100110101001101010001010011110101000101010001010100010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011011110110111111010100010110010111101001111101010110010,
	240'b101101001111111111101101101011101010011110101101110000001100110011001011110001111011110010110010101010101010100010101001101010101010101010101010101010101010101010101010101010101010100011011111111000001010100010110010111101001111101010110010,
	240'b101101001111111111101101101011001011100111101000111111011111111111111111111111111111110111110011111000111100110010110100101010011010100110101010101010101010101010101010101010101010100011010101110101101010100010110010111101001111101010110010,
	240'b101101001111111111101100101110001111000011111111111111111111111111111111111111111111111111111111111111111111111111110101110110001011010110101000101010011010101010101010101010101010101010101110101011101010100110110010111101001111101010110010,
	240'b101101001111111111101100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011001100101010111010100110101010101010101010101010101001101010011010100110110010111101001111101010110010,
	240'b101101001111111111110011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011011001010101000101010101010101010101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111111000111111001111111111111111111111111111111111111111111111111111111111111111111111111111101011110101111101101111111111111111111111111110101010110110101010001010101010101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111111000111111001111111111111111111111111111111111111111111111111111111111111111111111111101100110110011101101101101111111111111111111111111111111101101101101011010100010101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111110111111111001111111111111111111111111111111111111111111111111111111111111111111111111101001010100111101010001010111011100101111111111111111111111111111010011011000010101001101010101010100110110010111101001111101010110010,
	240'b101101001111111111110101111110101111111111111111111111111111111111111111111111111111111111111111111111111101001110101000101010101010011110110011111011111111111111111111111111111101101110101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111110010111100111111111111111111111111111111111111111111111111111111111111111111111111111101001110100111101100111011100110100111111000011111111111111111111111111111110111000110101010001010100110110010111101001111101010110010,
	240'b101101001111111111101110111010011111111111111111111111111111111111111111111111111111111111111111111111111101001110100110101110101110110010111000110111111111111111111111111111111111111111110000101100011010100010110010111101001111101010110010,
	240'b101101001111111111101011110110011111111111111111111111111111111111111111111111111111111111111111111111111101001110100110101110001111101111101101111010101111111111111111111111111111111111111111110100101010011010110010111101001111101010110010,
	240'b101101001111111111101011110001101111111011111111111111111111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111101111111111111111111111111111111111111111111100101011000010110001111101001111101010110010,
	240'b101101001111111111101100101101011111001011111111111111111111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111100100110110000111101001111101010110010,
	240'b101101001111111111101101101011001101101111111111111111111111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111110010010110011111101001111101010110010,
	240'b101101001111111111101101101010111011110111111100111111111111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111111011110111110111100111111101010110010,
	240'b101101001111111111101101101011011010101011100101111111111111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111111111011001111111100101111101010110010,
	240'b101101001111111111101101101011101010011110111111111111001111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111111111111100000111100111111100110110010,
	240'b101101001111111111101101101011101010100110101001110111001111111111111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111111111111101110111101001111100110110010,
	240'b101101001111111111101101101011101010100110101001101100101111000011111111111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111111111111110110111101101111100110110010,
	240'b101101001111111111101101101011101010100110101010101010001100000011111001111111111111111111111111111111111101001110100110101110001111100111111111111111111111111111111111111111111111111111111111111111111111111111111001111110011111100110110010,
	240'b101101001111111111101101101011101010100110101010101010101010100011001011111111001111111111111111111111111101001010100101101101111111100111111111111111111111111111111111111111111111111111111111111111111111111111111010111110101111100110110010,
	240'b101101001111111111101101101011101010100110101010101010101010101010101001110011011111110011111111111111111111000111100011111010001111110111111111111111111111111111111111111111111111111111111111111111111111111111111010111110101111100110110010,
	240'b101101001111111111101101101011101010100110101010101010101010101010101001101010011100100011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101111111100110110010,
	240'b101101001111111111101101101011101010100110101010101010101010101010101010101010101010100010111011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100111100111111100110110010,
	240'b101101001111111111101101101011101010100110101001101010011010101010101010101010101010101010101000101011101100110011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011000001111100111111101010110010,
	240'b101101001111111111101101101011011010101011010000110001011010100010101010101010101010101010101010101010011010100010110010110010101110100011111001111111111111111111111111111111111111111111111111111101011100001110110000111101001111101010110010,
	240'b101101001111111111101101101011011010101011101010110101111010011110101010101010101010101010101010101010101010101010101001101010001010110010111000110010001101011111100000111001001110010011010110101110001010011110110010111101001111101010110010,
	240'b101101001111111111101101101011011010101011101000110101101010011110101010101010101010101010101010101010101010101010101010101010101010100110101000101010001010100010101001101010101010101010101000101010011010100110110010111101001111101010110010,
	240'b101101001111111111101101101011011010101011101000110101101010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111101101101011011010100111101000110101101010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111101101101100001011000111100111110101101010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101001111101010110010,
	240'b101101001111111111101100101101101110000111110010110101001010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101001111101010110010,
	240'b101100011111111111110000101011111101110011111111110101001010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110011111101111111101010101111,
	240'b101001001111100111111100101111101010101111010000101111101010011110101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011011000110111111101111001110011101,
	240'b101101111101111011111111111100001100010010111000101110011011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101100100011110100111111111101011010110100,
	240'b111100011011100111110100111111111111111011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111011111100000111110100,
	240'b111111011101110010111011111001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100010101111001110110111111101,
	240'b111101001111111111101010101011001010000110101001101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101011101010111010101110101011101010011001111110101010111001011111001111110100,
	240'b111110011111011011100011100110011001001010101011101011011010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101010111001000010100100111011111111110011111001,
	240'b111111011110100010111100110010101110000011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001101111011001001110010101111101111111100,
	240'b111110101011110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011100101011111101,
	240'b110010111101000111111111111100111001100101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011011010111010001111111001111111111100110011001011,
	240'b101001001111010011111100011010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010110000000010000010111111111110110110011100,
	240'b101011101111111111011100000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110111100110100111100011111111011001111110010101011,
	240'b101101001111111111001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000111010001010111000100001110111001111110010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101001000011100000100011110111001111110010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101000000000000000011000110111101111110010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101000010000000000011000110111101111110010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101000010000000000011000110111101111110010110010,
	240'b101101001111111111001010000010110000000000001011010001000110011001100100010101110011011000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101001000000000000011000110111101111110010110010,
	240'b101101001111111111001010000001100010110110111011111110101111111111111111111111111111100011011100101011000110011100011111000000000000000000000000000000000000000000000000000000000000000010000011100001100000000000011000110111101111110010110010,
	240'b101101001111111111000101001010111101000111111111111111111111111111111111111111111111111111111111111111111111111111100000100010110010001100000000000000000000000000000000000000000000000000001100000011010000000000011001110111101111110010110010,
	240'b101101001111111111000110100110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101100111000001100000000000000000000000000000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111011011111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001000001100100000000000000000000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111101001111101101111111111111111111111111111111111111111111111111111111111111111111111111111000011100000111001011111111111111111111111111100000100100100000000000000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111101010111101101111111111111111111111111111111111111111111111111111111111111111111111111000111000011111001001101001111011111111111111111111111111001001001000110000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111100111111101011111111111111111111111111111111111111111111111111111111111111111111111110111101100000000000000000000111110110000111111111111111111111111101111010001001000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111100001111100011111111111111111111111111111111111111111111111111111111111111111111111110111110100000000000000000000000000011010110100001111111111111111111111111001010000000011000000000000000000011001110111101111110010110010,
	240'b101101001111111111010111110111001111111111111111111111111111111111111111111111111111111111111111111111110111110100000000000110110010111000000000101001001111111111111111111111111111100101010101000000000000000000011001110111101111110010110010,
	240'b101101001111111111001011101111001111111111111111111111111111111111111111111111111111111111111111111111110111110100000000001100001100011000101100101000001111111111111111111111111111111111010010000101100000000000011001110111101111110010110010,
	240'b101101001111111111000010100011001111111111111111111111111111111111111111111111111111111111111111111111110111110100000000001010111111010011001000101111111111111111111111111111111111111111111111011101110000000000011000110111101111110010110010,
	240'b101101001111111111000011010101001111101111111111111111111111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111011111111111111111111111111111111111111111110110100001001000010101110111101111110010110010,
	240'b101101001111111111000110001000011101100011111111111111111111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111110101111000010001110111101111110010110010,
	240'b101101001111111111001001000001111001010011111111111111111111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111111010111100011010110111011111110010110010,
	240'b101101001111111111001010000001010011100111110111111111111111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111111110011100111101110110011111110010110010,
	240'b101101001111111111001010000010100000010010110001111111111111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111111111110101110000110101101111110010110010,
	240'b101101001111111111001010000010110000000000111110111101011111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111111111111110100010110110001111110010110010,
	240'b101101001111111111001010000010110000000000000010100101011111111111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111111111111111001100110111011111101110110010,
	240'b101101001111111111001010000010110000000000000000000110101101001111111111111111111111111111111111111111110111110100000000001010111110110111111111111111111111111111111111111111111111111111111111111111111111111111100101111001001111101110110010,
	240'b101101001111111111001010000010110000000000000000000000000100001111101110111111111111111111111111111111110111110100000000001010101110110111111111111111111111111111111111111111111111111111111111111111111111111111101101111010111111101010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000001100100111101101111111111111111111111110111101100000000001010001110110111111111111111111111111111111111111111111111111111111111111111111111111111110000111011101111101010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000011010101111010111111111111111111101011010101011101110111111100111111111111111111111111111111111111111111111111111111111111111111111111111110001111011111111101010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000101101011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111001111111101010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000000000000110101101110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111110110101111110010110010,
	240'b101101001111111111001010000010110000000000000000000000000000000000000000000000000000000000000000000011000110011111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111110001101000101110110001111110010110010,
	240'b101101001111111111001010000010100000000001110010010100000000000000000000000000000000000000000000000000000000000000011000011000101011100111101100111111111111111111111111111111111111111111111111111000010100101000010011110111101111110010110010,
	240'b101101001111111111001010000010100000000010111111100001100000000000000000000000000000000000000000000000000000000000000000000000000000011000101011010110111000011010100011101100001011000010000100001010010000000000011000110111101111110010110010,
	240'b101101001111111111001010000010100000000010111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111001010000010100000000010111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111001010000010010000000010111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111001001000101000001011110110111100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001110111101111110010110010,
	240'b101101001111111111000110001001001010011011011000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110111011111110010110010,
	240'b101100011111111111010001000011111001010111111111011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111001001111110010101111,
	240'b101001001111101011110100001111000000011001110011001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111110111111010010011101,
	240'b101101111101111011111111110100010100111100101010001011100011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000101101111011110111111111101011010110100,
	240'b111100011011100111110101111111111111101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101111111011111111111011111100000111110100,
	240'b111111011101110010111011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100010101111001110110111111101,
	240'b111101001111111111101010101011001010000110101001101010101010101010101010101010101010101010101011101010111010101110101011101010101010101010101010101010101010101010101011101010111010101110101011101010011001111110101010111001011111001111110100,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule