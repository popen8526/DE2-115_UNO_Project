module wild_draw_four(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b110110011111111111011111100110101001110010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001001001010110111011111111011111111111111111,
	240'b110110111110110110111011110110011111001011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110100111001100110010011111110011111111,
	240'b110011111100001011110001111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111111111111111110101001101000111111010,
	240'b101010001110010011111111110111000110111001001111010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010010110100100101001110010011100100111001001110010101001001100111111010111111111100100011000001,
	240'b100110011111110111110001001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110100000100000000000000000000000000000000000000000000001010010111111111111101101110100101,
	240'b100101111111111111000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010101110000100100100000000000000000000000000000000000000000001000010111111001110111010111000,
	240'b100110011111111110110001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100010001111111000000000000000000000000000000000000000000110111111101111111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011100011001000010011010001000100100000000000001110100101010001010100110001111101111111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111001100100010011001110010111110001001001101100111110010111001101010010111101001111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100111001000011100010001001101110100100100111110100111111101111010010001111111011111111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110111111111011110110011110001111011100010000000111010111101000100100000111110111101101111001010111101,
	240'b100110101111111110110010000000010000000000100110011100011001010010001101011110110101011100110001000011010000000000000000000000000000000101101001111101101000010101100100010110010000100000001000010111100000110100110100111101111111001010111101,
	240'b100110101111111110110001000000000101111011100100111111111111111111111111111111111111111111110110110011011000101000110100000000010000000000011000101000010001110000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110101100010010011111001011111111111111111111111111111101111010001110010011100101111010011110100111011001101000000011011000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110111000101111101111111111111111111111111111111111001111110000001101010111010111110101101101011111010010110100001110101001111111000010110000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111010111111100011111111111111111111111111111111111001010111100101101010110100010101000011010010111011100110110111110000111111111101100010010000100000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111101000111110001111111111111111111111111111111111100010110110111001000001001011010100000100111001101110110111001100111011111111111111111100111100101011000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111101000111101111111111111110011111010101110101111011100110000011001100101001010010101010101010001010011110001011100011011100110111010111111010011001111001001110000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111100010111101111111000110110011110010101100111111001111110001111100010110001110010100100101010101010000101001001100010110111010110010111100011011011010101111110001001100000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111010111111101001110100111010001111101101011010110101001101010101100101111110110011100000101000101010001011111111101100111011111111111111111111111001110111100101001010100000010000000000000000000111000111101111111001010111101,
	240'b100110011111111111001000111000111111100111001101110001010101001001010000010100000101010111001001100111010100110101010011011000111101011111001110111111111111111111100000110110111111101001001111000000000000000000111000111101111111001010111101,
	240'b100110101111111110111000110000011111111111001100110100100101110001010011010101010100111110010100110001000100101101001101010011001011110111001101111110101111111111110100110010001111111111001010000011110000000000111000111101111111001010111101,
	240'b100110101111111110101011100100101111111111011000110110010111011001010001010101010101001001110010110101111001010110101010101001111011000011000100111011011111111111111101110010001111100011111111011001110000000000111000111101111111001010111101,
	240'b100110101111111110101011010101011111111011101010110101011001100001010000010101010101010001011010110100011101000011111111111111111110100010110010110111001111111111111111110011111110101011111111110010100000100000110101111101111111001010111101,
	240'b100110101111111110101111000111001110000011111011110011001011110001010010010101010101010101010001101100111100111111110100111111111111110010110111110010101111111111111111111000111101010111111111111111000100010100110000111101111111001010111101,
	240'b100110101111111110110010000000001001100111111111110011011101001101011111010100110101010101010000100100001101010111100101111111111111111110111111101101011111111011111111111100111100101011111111111111111001010000110011111101101111001010111101,
	240'b100110011111111110110010000000000011110011111001110110111101101001111000010100010101010101010010011011101101101011010011111111111111111111001111110011101111111111111111111111111100011011111000111111111101001101001010111101001111001010111101,
	240'b100110011111111110110010000000010000010010110001111100011101001110011101010011000101001001010001010101101100110111001101111111011111111111101100110100001111111111111111111111111101001111100111111111111111000101110010111100001111001010111101,
	240'b100110011111111110110010000000100000000000111110111100001100101111011111100000000110111001101111011101111110001111001100111101001111111111111001110001111111111011111111111111111110010111010110111111111111111110011111111011111111001010111101,
	240'b100110011111111110110010000000100000000000000001100011111101011111011111111001011101110011011101111000011110111011000000111011011111111111111111110010011110001011101101111011011101110111000111111111111111111111000110111100011111001010111101,
	240'b100110011111111110110010000000100000000000000000000101101100010111011000110010011100101110101111101111011100011111010000111111011111111111111111110101101010111111001001110010001100011011101101111111111111111111100100111100111111000110111101,
	240'b100110011111111110110010000000100000000000000000000000000011010011100111111111111111111111011100111000101111111111111111111111111111111111111111111011001101000111111111111111111111111111111111111111111111111111101101111101001111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000001001011111011001111111111101111110011001111111111111111111111111111111111111111111111001100011111111100111111111111111111111111111111111111111111110000111101101111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000010011101110010011111111110010001110011011110001111100011111000111110001111011111011111011110101111111111111111111111111111111111111111111110000111101011111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000011100111001110111110001100111011001101110011101100111011001110110010011101010011111110111111111111111111111111111111111111111111010110111100101111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000000000011000100100111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000100111100001111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000101100001001000000000100000010101101111100111111111111111111111111111111111111111111111111111111111111111111111111111001101100111100111101011111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000111110010010010000000000000000000000101001101111000010011000010111010111111100011111111111111111111111111110010100110110001000000110100111101111111001010111101,
	240'b100110011111111110110010000000000101000101011001000000000100001010010011100101011101011111100010001110010000000000000000000000000000000000001010001000110100011001011111011010110110010100110110000000100000000000111000111101111111001010111101,
	240'b100110011111111110110011001011101011100011000010001011000111011011111111110010111110100111101111010011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111110111000101110001111110111111101101110100011111111011111001010111000111110101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111110110011001001001011001010111101001001000000010010110010100010111001001110110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110110010000000000100100001001111000000000000000001010000110110100110010001001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000001011110010100111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111101111111001010111101,
	240'b100110011111111111000111000001110000000000000000000000000000000000000000011010111100101000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001111111011110110010110110,
	240'b100110111111101111110111010101010000000000000000000000000000000000000000000001000011000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110101010111111111101100010100110,
	240'b101011101101110111111111111010111001010001111000011110100111101001111010011110000111010001111001011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111001011111011011100011111111111111001100011011001101,
	240'b110011111100000011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010101101001111111001,
	240'b110011011110100011000000110011001110010111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100001101101010111111110010011111000011110000,
	240'b110010111111011011100011101001101010101010110101101101101011010110110101101101011011010110110101101101101011011010110110101101101011011010110101101101011011010110110101101101101011011010110110101100101010001110110010111011001111000011101111,
	240'b110110011111111111011111100110101001110010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001001001010110111011111111011111111111111111,
	240'b110110111110110110111011110110011111001011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110100111001100110010011111110011111111,
	240'b110011111100001011110001111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111111111111111110101001101000111111010,
	240'b101010001110010011111111110111000110111001001111010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010010110100100101001110010011100100111001001110010101001001100111111010111111111100100011000001,
	240'b100110011111110111110001001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110100000100000000000000000000000000000000000000000000001010010111111111111101101110100101,
	240'b100101111111111111000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010101110000100100100000000000000000000000000000000000000000001000010111111001110111010111000,
	240'b100110011111111110110001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100010001111111000000000000000000000000000000000000000000110111111101111111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011100011001000010011010001000100100000000000001110100101010001010100110001111101111111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111001100100010011001110010111110001001001101100111110010111001101010010111101001111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100111001000011100010001001101110100100100111110100111111101111010010001111111011111111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110111111111011110110011110001111011100010000000111010111101000100100000111110111101101111001010111101,
	240'b100110101111111110110010000000010000000000100110011100011001010010001101011110110101011100110001000011010000000000000000000000000000000101101001111101101000010101100100010110010000100000001000010111100000110100110100111101111111001010111101,
	240'b100110101111111110110001000000000101111011100100111111111111111111111111111111111111111111110110110011011000101000110100000000010000000000011000101000010001110000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110101100010010011111001011111111111111111111111111111101111010001110010011100101111010011110100111011001101000000011011000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110111000101111101111111111111111111111111111111111001111110000001101010111010111110101101101011111010010110100001110101001111111000010110000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111010111111100011111111111111111111111111111111111001010111100101101010110100010101000011010010111011100110110111110000111111111101100010010000100000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111101000111110001111111111111111111111111111111111100010110110111001000001001011010100000100111001101110110111001100111011111111111111111100111100101011000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111101000111101111111111111110011111010101110101111011011110000011001100101001010010101010101010001010011110001011100011011100110111010111111010011001111001001110000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111100010111101111111000110110011110010011100110111001100110001011100001110001110010100100101010101010000101001001100010110111101110100001100100011011010101111110001001100000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111010111111101001110100111010000111111011101110011010110110101111110100011111000011011110101000101010001100000001101011110011010101101001110110111010000111100101001010100000010000000000000000000111000111101111111001010111101,
	240'b100110011111111111001000111000111111100111001011111000101010100010101000101010001010101011100111100110110100110101010011011000111101100101101000010010111000100011011100110111001111101001001111000000000000000000111000111101111111001010111101,
	240'b100110101111111110111000110000011111111111001010111000111010111010101001101010101010011111001100110000110100101101001101010011001100001110001110010011000101111111010101110011001111111111001010000011110000000000111000111101111111001010111101,
	240'b100110101111111110101011100100101111111111010111110111101011110010101000101010101010100010111010110111101001010110101101101010011011001110101001010011100101001110111101110011011111100011111111011001110000000000111000111101111111001010111101,
	240'b100110101111111110101011010101011111111011101001110100111100110110100111101010101010100110101101111001011011110011011101111101001110101010101100010110000100111110011011110100111110101011111111110010100000100000110101111101111111001010111101,
	240'b100110101111111110101111000111001110000011111011110010011101110110101001101010101010101010101000110110111011010010011110101100101110101110111101011010000100111001110111110110111101011111111111111111000100010100110000111101111111001010111101,
	240'b100110101111111110110010000000001001100111111111110010111110001110110000101010011010101010100111110010101100110010011010101010001101100111000101011000100101000001011110110100101100111011111111111111111001010000110011111101101111001010111101,
	240'b100110011111111110110010000000000011110011111001110110101101111010111101101010001010101010101000101110001110000110010111101010001100100011001000010011010101010001010010101110111100101111111001111111111101001101001010111101001111001010111101,
	240'b100110011111111110110010000000010000010010110001111100011101001011010000101001101010100010101000101010111110010110100010101001101011011011100011011000000101000001001100100101101101010111100111111111111111000101110010111100001111001010111101,
	240'b100110011111111110110010000000100000000000111110111100001100101011101111110000011011100010111000101111001111010110110110101000001010110011100110100010100110101001101101101011111110011011010110111111111111111110011111111011111111001010111101,
	240'b100110011111111110110010000000100000000000000001100011111101011111011110111010101110010111100101111010001110111110110001100111011010100111010111110001111101000111011101111010101101111011000111111111111111111111000110111100011111001010111101,
	240'b100110011111111110110010000000100000000000000000000101101100010111011000110010001100101010101110101101111001110010010010101010001010100011000101110101011011001011001011110010001100010111101101111111111111111111100100111100111111000110111101,
	240'b100110011111111110110010000000100000000000000000000000000011010011100111111111111111111111011100110111111100001010101000101010011010100010110011111000101101001111111111111111111111111111111111111111111111111111101101111101001111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000001001011111011001111111111101111110011011110100010111000101101001011010010111111111101001100100011111100111111111111111111111111111111111111111111110000111101101111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000010011101110010011111111110010001110011111101010111001111110011111101011111011111011111011110101111111111111111111111111111111111111111111110000111101011111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000011100111001110111110001100111011001110110011111100111111001111110010011101010011111110111111111111111111111111111111111111111111010110111100101111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000000000011000100100111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000100111100001111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000101100001001000000000100000010101101111100111111111111111111111111111111111111111111111111111111111111111111111111111001101100111100111101011111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000111110010010010000000000000000000000101001101111000010011000010111010111111100011111111111111111111111111110010100110110001000000110100111101111111001010111101,
	240'b100110011111111110110010000000000101000101011001000000000100001010010011100101011101011111100010001110010000000000000000000000000000000000001010001000110100011001011111011010110110010100110110000000100000000000111000111101111111001010111101,
	240'b100110011111111110110011001011101011100011000010001011000111011011111111110010111110100111101111010011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111110111000101110001111110111111101101110100011111111011111001010111000111110101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111110110011001001001011001010111101001001000000010010110010100010111001001110110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110110010000000000100100001001111000000000000000001010000110110100110010001001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000001011110010100111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111101111111001010111101,
	240'b100110011111111111000111000001110000000000000000000000000000000000000000011010111100101000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001111111011110110010110110,
	240'b100110111111101111110111010101010000000000000000000000000000000000000000000001000011000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110101010111111111101100010100110,
	240'b101011101101110111111111111010111001010001111000011110100111101001111010011110000111010001111001011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111001011111011011100011111111111111001100011011001101,
	240'b110011111100000011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010101101001111111001,
	240'b110011011110100011000000110011001110010111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100001101101010111111110010011111000011110000,
	240'b110010111111011011100011101001101010101010110101101101101011010110110101101101011011010110110101101101101011011010110110101101101011011010110101101101011011010110110101101101101011011010110110101100101010001110110010111011001111000011101111,
	240'b110110011111111111011111100110101001110010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001001001010110111011111111011111111111111111,
	240'b110110111110110110111011110110011111001011111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110100111001100110010011111110011111111,
	240'b110011111100001011110001111111111111111111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111111111111111111110101001101000111111010,
	240'b101010001110010011111111110111000110111001001111010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010010110100100101001110010011100100111001001110010101001001100111111010111111111100100011000001,
	240'b100110011111110111110001001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110100000100000000000000000000000000000000000000000000001010010111111111111101101110100101,
	240'b100101111111111111000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010101110000100100100000000000000000000000000000000000000000001000010111111001110111010111000,
	240'b100110011111111110110001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100010001111111000000000000000000000000000000000000000000110111111101111111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011100011001000010011010001000100100000000000001110100101010001010100110001111101111111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111001100100010011001110010111110001001001101100111110010111001101010010111101001111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100111001000011100010001001101110100100100111110100111111101111010010001111111011111111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110111111111011110110011110001111011100010000000111010111101000100100000111110111101101111001010111101,
	240'b100110101111111110110010000000010000000000100110011100011001010010001101011110110101011100110001000011010000000000000000000000000000000101101001111101101000010101100100010110010000100000001000010111100000110100110100111101111111001010111101,
	240'b100110101111111110110001000000000101111011100100111111111111111111111111111111111111111111110110110011011000101000110100000000010000000000011000101000010001110000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110101100010010011111001011111111111111111111111111111101111010001110010011100101111010011110100111011001101000000011011000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110111000101111101111111111111111111111111111111111001111110000001101001011010010110100101101001011001111110100001110101001111111000010110000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111010111111100011111111111111111111111111111111111001010111100001111111111111111111111111111111111111111110110101110000111111111101100010010000100000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111101000111110001111111111111111111111111111111111100001110110111111111111111111111111111111111111111111111011111100110011111111111111111100111100101011000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111101000111101111111111111110011111010101110101111011011101111011110101111110101111111111111111111111111111111001100000111100110111010111111010011001111001001110000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111100010111101111111000110110011110010101100111111001111110001101100110111000101111010101111111111111111111111111100000010111101110100001100100011011010101111110001001100000000000000000000000000111000111101111111001010111101,
	240'b100110011111111111010111111101001110100111010001111101101011010110101001101010101100101011101111110010011111111011111111111111111101110010011001101101001110110111010000111100101001010100000010000000000000000000111000111101111111001010111101,
	240'b100110011111111111001000111000111111100111001101110001010101001001010000010100000101010111000100110010111111011111111111111111111111001101100101010010111000100011011100110111001111101001001111000000000000000000111000111101111111001010111101,
	240'b100110101111111110111000110000011111111111001100110100100101110001010011010101010100111110010001110101111101100011101110111011101111101110001001010011000101111111010101110011001111111111001010000011110000000000111000111101111111001010111101,
	240'b100110101111111110101011100100101111111111011000110110010111011001010001010101010101001001110010110101111010110111001110110011001100110010101000010011100101001110111101110011011111100011111111011001110000000000111000111101111111001010111101,
	240'b100110101111111110101011010101011111111011101010110101011001100001010000010101010101010001011010110101001001100110001011110010011110100110101100010110000100111110011011110100111110101011111111110010100000100000110101111101111111001010111101,
	240'b100110101111111110101111000111001110000011111011110011001011110001010010010101010101010101010001101110101000011100000000000101001100100011000000011010000100111001110111110110111101011111111111111111000100010100110000111101111111001010111101,
	240'b100110101111111110110010000000001001100111111111110011011101001101011111010100110101010101010000100101001011110000000100000000001000011011001010011000100101000001011110110100101100111011111111111111111001010000110011111101101111001010111101,
	240'b100110011111111110110010000000000011110011111001110110111101101001111000010100010101010101010010011011111101101000100011000000000100111111001000010011100101010001010010101110111100101111111001111111111101001101001010111101001111001010111101,
	240'b100110011111111110110010000000010000010010110001111100011101001110011101010011000101001001010001010101101101010001010100000000000010000011010001011000100101000001001100100101101101010111100111111111111111000101110010111100001111001010111101,
	240'b100110011111111110110010000000100000000000111110111100001100101111011111100000000110111001101111011101111110100110001110000000000000001110110110100011100110101001101101101011111110011011010110111111111111111110011111111011111111001010111101,
	240'b100110011111111110110010000000100000000000000001100011111101011111011111111001011101110011011100111000011111001110010100000000000000000010000001110011001101000111011101111010101101111011000111111111111111111111000110111100011111001010111101,
	240'b100110011111111110110010000000100000000000000000000101101100010111011000110010011100101110110001101011000100010100010111000000000000000001001010110100111011001111001011110010001100010111101101111111111111111111100100111100111111000110111101,
	240'b100110011111111110110010000000100000000000000000000000000011010011100111111111111111111111011101110110100011101000000000000000000000000000010111110011111101010111111111111111111111111111111111111111111111111111101101111101001111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000001001011111011001111111111101111110100011011001000101010000111000001101100111011111000101100101011111100111111111111111111111111111111111111111111110000111101101111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000010011101110010011111111110010001110100011011011110100101101000111011110111011111011111011110101111111111111111111111111111111111111111111110000111101011111000110111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000011100111001110111110001100111011010001110100101101001011010001110010011101010011111110111111111111111111111111111111111111111111010110111100101111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000000000011000100100111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000100111100001111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000000000000000000000101100001001000000000100000010101101111100111111111111111111111111111111111111111111111111111111111111111111111111111001101100111100111101011111001010111101,
	240'b100110011111111110110010000000100000000000000000000000000000000000000000000000000111110010010010000000000000000000000101001101111000010011000010111010111111100011111111111111111111111111110010100110110001000000110100111101111111001010111101,
	240'b100110011111111110110010000000000101000101011001000000000100001010010011100101011101011111100010001110010000000000000000000000000000000000001010001000110100011001011111011010110110010100110110000000100000000000111000111101111111001010111101,
	240'b100110011111111110110011001011101011100011000010001011000111011011111111110010111110100111101111010011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111110111000101110001111110111111101101110100011111111011111001010111000111110101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110011111111110110011001001001011001010111101001001000000010010110010100010111001001110110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110110010000000000100100001001111000000000000000001010000110110100110010001001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111101111111001010111101,
	240'b100110101111111110110010000000100000000000000000000000000000000000001011110010100111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111101111111001010111101,
	240'b100110011111111111000111000001110000000000000000000000000000000000000000011010111100101000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001111111011110110010110110,
	240'b100110111111101111110111010101010000000000000000000000000000000000000000000001000011000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110101010111111111101100010100110,
	240'b101011101101110111111111111010111001010001111000011110100111101001111010011110000111010001111001011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111001011111011011100011111111111111001100011011001101,
	240'b110011111100000011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010101101001111111001,
	240'b110011011110100011000000110011001110010111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100001101101010111111110010011111000011110000,
	240'b110010111111011011100011101001101010101010110101101101101011010110110101101101011011010110110101101101101011011010110110101101101011011010110101101101011011010110110101101101101011011010110110101100101010001110110010111011001111000011101111,
};
assign data = picture[addr];
endmodule