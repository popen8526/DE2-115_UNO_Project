module red_skip(
    input [7:0] addr,
    output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100001111001111110010110011101011010110110110101101111011011010110110101101101011011010110110101101111011011110110111101101111011011010110110101101101011011010110110101101101011011110110111101101101011010111000110111010011111001011110000,
	240'b111100011110100011000000110100101111000011110011111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100111111001011010101101110001110000111110001,
	240'b111011011011110011100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011100111101010,
	240'b101110001101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010111000,
	240'b100110111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010011111,
	240'b101011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101101101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111000,
	240'b101100101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011,
	240'b100111111111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110100010,
	240'b101010101101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110101011,
	240'b111001001011101011110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011011110011100000,
	240'b111100101101101110111101111010111111111111111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111111101111101111011101001011110010,
	240'b111110011111110011100011101000111001011110101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001001101110011111111000011111110011111001,
	240'b111100001111001111110011110011101011011010110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011010111000110111010101111001111110000,
	240'b111100011110100011000000110100101111000011110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001011010101101110001110000111110001,
	240'b111011011011110011100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011100111101010,
	240'b101110001101000011111111111101001011000010001100100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010100001111000011010001000100010101010100011101110111111111101101010111000,
	240'b100110111111000011111110100111010100111101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100111001010101011110011000100101101100010011110100110110001100111110101111101010011111,
	240'b101011111111111011101110011001100101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110011011001000111100111111000011110010101010000101010001011100111000001111111110101111,
	240'b101101101111111111100101011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101011100000011111111101100100110110010100010111101101001001001010101110101101111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011100101110110111011011111001110111001101001010101101011101011001011101110101011111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100010111110010001101111110011101110010101100111100001011110010101101011110101001111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000111110101101100111011000011101110011010011101001101110000101100110110101001111111110111000,
	240'b101101101111111111100101011000100101001101010011010100000101000101010001010100000101000001010010010101000101010101010101010101010101010101010011011000111110011110110001010100000110101111100011111111011011101001011000110101101111111110111000,
	240'b101101011111111111100101011000100100111101011110100010101010001010100010100110101000100101110011010111000101001001010001010101000101010101010101010100011001001111110110110011011011000011101011111001100110111001010111110101101111111110111000,
	240'b101101011111111111100101010111100111001011010100111111101111111111111111111111111111111011110010110110101010111101111011010101100101000101010100010101010101010010001010110011111101111010111101011100010101000101011010110101101111111110111000,
	240'b101101011111111111100011011101001101111111111111111111111111111111111111111111111111111111111111111111111111111111110110110001100111111001010011010100110101010101010001010110000101110101010100010100100101010001011010110101101111111110111000,
	240'b101101011111111111100010101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110110011011000110101000101010101010101000101001101010100010101010101010001011010110101101111111110111000,
	240'b101101011111111111101100111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111011001010000010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101101011111111111110011111110011111111111111111111111111111111111111111111111111111111111111111111111111111100011101110111011011111011111111111111111111110101010000001010100000101010101010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111110100111110011111111111111111111111111111111111111111111111111111111111101011101010110111100101100101011001000111011010100011111000111111111111101101011111010101000001010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111110010111110011111111111111111111111111111111111111111111111111100111001101110010100000100111001001101010011010100111001001111011001111100000111111111111001110110111001010001010101010101010001011010110101101111111110111000,
	240'b101101101111111111101111111100111111111111111111111111111111111111111111110100100110000001010000010101100110101110000110100001100110111001010011010011110101100111000010111111111101000001011100010100110101010001011010110101101111111110111000,
	240'b101101101111111111101001111000011111111111111111111111111111111111110000011101000101000001010010011011101110001111111111111111111110111010101110010111010100111101100111111001011111111110100110010100010101010001011010110101101111111110111000,
	240'b101101101111111111100011110010111111111111111111111111111111111110110010010100010101001101010010010101101010011011111110111111111111111111111111101111000101011101001110100111111111111111110001011100110101000001011010110101101111111110111000,
	240'b101101011111111111100000101010011111111111111111111111111111100101111100010011100111000001101110010100000101010110110010111111111111111111111111111111011000101101001101011011011111000111111111101111010101001001011010110101101111111110111000,
	240'b101101011111111111100001100001101111011111111111111111111110011101100010010011111011010111011011011001100100111101011001110000001111111111111111111111111100010101010010010110001101100011111111111101000111001001010110110101101111111110111000,
	240'b101101011111111111100100011010011101101011111111111111111101101001010111010100111101000111111111110010110101111001001111011000001100110111111111111111111101111101011100010100101100011011111111111111111010110101010110110101101111111110111000,
	240'b101101011111111111100101010111011010100111111111111111111101011101010110010101001101010111111111111111111011111001011001010011110110011111011001111111111110001001011110010100101100010011111111111111111101111101100100110101011111111110111000,
	240'b101101011111111111100101010111100111000011110011111111111110001001011101010100011011111011111111111111111111111110110000010101010100111101110000111010001101001101010101010101011101001011111111111111111111101110000101110100101111111110111000,
	240'b101101011111111111100101011000010101001010111110111111111111010001110010010011011000110011111110111111111111111111111101101000100101001001001111011111111000111101010000011001011110101011111111111111111111111110101101110100011111111110111000,
	240'b101101101111111111100101011000100100111101110100111100111111111110100000010011100101101011001001111111111111111111111111111110011001010101010011010100110101010001001111100011011111110111111111111111111111111111001101110101101111111110111000,
	240'b101101101111111111100101011000100101001101010010101011001111111111100010011000110100111101100110110010011111110111111111111111111111010001111010010100100101001101011010110100111111111111111111111111111111111111100110110111101111111110111000,
	240'b101101101111111111100101011000100101001101010011010111111101100011111111101101010101010001010000010111001000101110110000101100011001001001100001010100100101000110100101111111101111111111111111111111111111111111110010111001101111111110111000,
	240'b101101101111111111100101011000100101001101010101010100010111011111101101111111101010100101011000010011110100111101010001010100010100111101001111010101011001110011111000111111111111111111111111111111111111111111110110111011011111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101000010001010111101001111111111001001100000000101110001010101010101010101101101111010110000001111110011111111111111111111111111111111111111111111111111111000111100011111111110111000,
	240'b101101011111111111100101011000100101001101010101010101010101010101010001100011111111010011111111111110001101111011000111110001111101101111110110111111111111111111111111111111111111111111111111111111111111111111111000111100101111111110111000,
	240'b101101011111111111100101011000100101001101010101010101010101010101010100010100011000011011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111010011111111110111000,
	240'b101101011111111111100101011000100101001101010101010101010101010101010101010101010101000001110010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110110011111111110111000,
	240'b101101011111111111100101011000100101001101010100010100010101001001010001010100100101010101010001010110101001011011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001110110100101111111110111000,
	240'b101101011111111111100101011000100101000101011000100010111011001110101000011100010101001001010101010101000101000001100011100101111101000111110100111111111111111111111111111111111111111111111111111101101001111101011001110101101111111110111000,
	240'b101101011111111111100101011000000101011110111001111101101110000011101011111011101000010101010001010101010101010101010011010100000101100101110001100101011011000011000100110011111101000110111001011111100101001001011001110101101111111110111000,
	240'b101101101111111111100101010111011001001011111111111010000110110101011111110000011110010101100011010100110101010101010101010101010101010001010010010100000101000001010110010110010101100101010011010100010101010001011010110101101111111110111000,
	240'b101101101111111111100101011000011100110111001011111000001100101101011000011001011110101110001101010100000101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111100100011001111101110110010110011100111111000010111110010110101101110110100000010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111100101011000011101000010110110010010101000010011110010101111101110100110001110010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111100101010111011001011111110011100001110101010110100000111111111110010101100100010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101100101111111111101010011000010101100010111111111101101101100111100100111011101000100001010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110101111111110110011,
	240'b100111111111011011111011100001010100101101011000100011011011011110101010011100100101000001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100111001110101111101001111111010100010,
	240'b101010101101110011111111111000011000010101101000011001100110011001100110011001110110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010010111110111010110111111111110011010101011,
	240'b111001001011101011110100111111111111101011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111100011111111111110011011110011100000,
	240'b111100101101101110111101111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111011101001011110010,
	240'b111110011111110011100011101000111001011110101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001001101110011111111000011111110011111001,
	240'b111100001111001111110010110011101011010110110110101101111011011010110110101101101011011010110110101101111011011110110111101101111011011010110110101101101011011010110110101101101011011110110111101101101011010111000110111010011111001011110000,
	240'b111100011110100011000000110100101111000011110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001011010101101110001110000111110001,
	240'b111011011011110011100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001011100111101010,
	240'b101110001101000011111111111101001011000010001100100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001010100001111000011010001000100010101010100011101110111111111101101010111000,
	240'b100110111111000011111110100111010100111101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010100111001010101011110011000100101101100010011110100110110001100111110101111101010011111,
	240'b101011111111111011101110011001100101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110011011001000111100111111000011110010101010000101010001011100111000001111111110101111,
	240'b101101101111111111100101011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101011100000011111111101100100110110010100010111101101001001001010101110101101111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011100101110110111011011111001110111001101001010101101011101011001011101110101011111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100010111110010001101111110011101110010101100111100001011110010101101011110101001111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100000111110101101100111011000011101110011010011101001101110000101100110110101001111111110111000,
	240'b101101101111111111100101011000100101001101010011010100000101000101010001010100000101000001010010010101000101010101010101010101010101010101010011011000111110011110110001010100000110101111100011111111011011101001011000110101101111111110111000,
	240'b101101011111111111100101011000100100111101011110100010101010001010100010100110101000100101110011010111000101001001010001010101000101010101010101010100011001001111110110110011011011000011101011111001100110111001010111110101101111111110111000,
	240'b101101011111111111100101010111100111001011010100111111101111111111111111111111111111111011110010110110101010111101111011010101100101000101010100010101010101010010001010110011111101111010111101011100010101000101011010110101101111111110111000,
	240'b101101011111111111100011011101001101111111111111111111111111111111111111111111111111111111111111111111111111111111110110110001100111111001010011010100110101010101010001010110000101110101010100010100100101010001011010110101101111111110111000,
	240'b101101011111111111100010101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110110011011000110101000101010101010101000101001101010100010101010101010001011010110101101111111110111000,
	240'b101101011111111111101100111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111011001010000010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101101011111111111110011111110011111111111111111111111111111111111111111111111111111111111111111111111111111100011101110111011011111011111111111111111111110101010000001010100000101010101010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111110100111110011111111111111111111111111111111111111111111111111111111111101011101010110111100101100101011001000111011010100011111000111111111111101101011111010101000001010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111110010111110011111111111111111111111111111111111111111111111111100111001101110010100000100111001001101010011010100111001001111011001111100000111111111111001110110111001010001010101010101010001011010110101101111111110111000,
	240'b101101101111111111101111111100111111111111111111111111111111111111111111110100100110000001010000010101100110101110000110100001100110111001010011010011110101100111000010111111111101000001011100010100110101010001011010110101101111111110111000,
	240'b101101101111111111101001111000011111111111111111111111111111111111110000011101000101000001010010011011101110001111111111111111111110111010101110010111010100111101100111111001011111111110100110010100010101010001011010110101101111111110111000,
	240'b101101101111111111100011110010111111111111111111111111111111111110110010010100010101001101010010010101101010011011111110111111111111111111111111101111000101011101001110100111111111111111110001011100110101000001011010110101101111111110111000,
	240'b101101011111111111100000101010011111111111111111111111111111100101111100010011100111000001101110010100000101010110110010111111111111111111111111111111011000101101001101011011011111000111111111101111010101001001011010110101101111111110111000,
	240'b101101011111111111100001100001101111011111111111111111111110011101100010010011111011010111011011011001100100111101011001110000001111111111111111111111111100010101010010010110001101100011111111111101000111001001010110110101101111111110111000,
	240'b101101011111111111100100011010011101101011111111111111111101101001010111010100111101000111111111110010110101111001001111011000001100110111111111111111111101111101011100010100101100011011111111111111111010110101010110110101101111111110111000,
	240'b101101011111111111100101010111011010100111111111111111111101011101010110010101001101010111111111111111111011111001011001010011110110011111011001111111111110001001011110010100101100010011111111111111111101111101100100110101011111111110111000,
	240'b101101011111111111100101010111100111000011110011111111111110001001011101010100011011111011111111111111111111111110110000010101010100111101110000111010001101001101010101010101011101001011111111111111111111101110000101110100101111111110111000,
	240'b101101011111111111100101011000010101001010111110111111111111010001110010010011011000110011111110111111111111111111111101101000100101001001001111011111111000111101010000011001011110101011111111111111111111111110101101110100011111111110111000,
	240'b101101101111111111100101011000100100111101110100111100111111111110100000010011100101101011001001111111111111111111111111111110011001010101010011010100110101010001001111100011011111110111111111111111111111111111001101110101101111111110111000,
	240'b101101101111111111100101011000100101001101010010101011001111111111100010011000110100111101100110110010011111110111111111111111111111010001111010010100100101001101011010110100111111111111111111111111111111111111100110110111101111111110111000,
	240'b101101101111111111100101011000100101001101010011010111111101100011111111101101010101010001010000010111001000101110110000101100011001001001100001010100100101000110100101111111101111111111111111111111111111111111110010111001101111111110111000,
	240'b101101101111111111100101011000100101001101010101010100010111011111101101111111101010100101011000010011110100111101010001010100010100111101001111010101011001110011111000111111111111111111111111111111111111111111110110111011011111111110111000,
	240'b101101101111111111100101011000100101001101010101010101010101000010001010111101001111111111001001100000000101110001010101010101010101101101111010110000001111110011111111111111111111111111111111111111111111111111111000111100011111111110111000,
	240'b101101011111111111100101011000100101001101010101010101010101010101010001100011111111010011111111111110001101111011000111110001111101101111110110111111111111111111111111111111111111111111111111111111111111111111111000111100101111111110111000,
	240'b101101011111111111100101011000100101001101010101010101010101010101010100010100011000011011101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111010011111111110111000,
	240'b101101011111111111100101011000100101001101010101010101010101010101010101010101010101000001110010110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110110011111111110111000,
	240'b101101011111111111100101011000100101001101010100010100010101001001010001010100100101010101010001010110101001011011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001110110100101111111110111000,
	240'b101101011111111111100101011000100101000101011000100010111011001110101000011100010101001001010101010101000101000001100011100101111101000111110100111111111111111111111111111111111111111111111111111101101001111101011001110101101111111110111000,
	240'b101101011111111111100101011000000101011110111001111101101110000011101011111011101000010101010001010101010101010101010011010100000101100101110001100101011011000011000100110011111101000110111001011111100101001001011001110101101111111110111000,
	240'b101101101111111111100101010111011001001011111111111010000110110101011111110000011110010101100011010100110101010101010101010101010101010001010010010100000101000001010110010110010101100101010011010100010101010001011010110101101111111110111000,
	240'b101101101111111111100101011000011100110111001011111000001100101101011000011001011110101110001101010100000101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111100100011001111101110110010110011100111111000010111110010110101101110110100000010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111100101011000011101000010110110010010101000010011110010101111101110100110001110010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101101101111111111100101010111011001011111110011100001110101010110100000111111111110010101100100010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110101101111111110111000,
	240'b101100101111111111101010011000010101100010111111111101101101100111100100111011101000100001010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011011110110101111111110110011,
	240'b100111111111011011111011100001010100101101011000100011011011011110101010011100100101000001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100111001110101111101001111111010100010,
	240'b101010101101110011111111111000011000010101101000011001100110011001100110011001110110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010010111110111010110111111111110011010101011,
	240'b111001001011101011110100111111111111101011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111100011111111111110011011110011100000,
	240'b111100101101101110111101111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111011101001011110010,
	240'b111110011111110011100011101000111001011110101111101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001001101110011111111000011111110011111001,
};
assign data = picture[addr];
endmodule