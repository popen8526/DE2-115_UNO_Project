module yellow_six(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111101111111100011101101101100111010010010111001101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101101101010001110111111111100101111011111110111,
	240'b111111111111111111011001101101101011110111010101110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110100101011101111000000111011111111111111111101,
	240'b111111101110100010111101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101111111111010011110100,
	240'b110100011100010111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001100101011000111,
	240'b101010011100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011110111100,
	240'b101011111101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001011000101,
	240'b101111101110001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111001011,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001101,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111001100,
	240'b101110011101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111011001001,
	240'b101001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100111000000,
	240'b101100101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011101110111010,
	240'b111010101101000011011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001101110011011100,
	240'b111111101111011110111101110101101111101011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111011011001110110010101111110111111011,
	240'b111100011111010111111001110000001010000010101000101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101011101010111010101110101011101001111001111011000001111100101111000111110011,
	240'b111101111111100011101101101100111010010010111001101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101101101010001110111111111100101111011111110111,
	240'b111111111111111111011001101101101011110111010101110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110100101011101111000000111011111111111111111101,
	240'b111111101110100010111101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101111111111010011110100,
	240'b110100011100010111110010111111111111001111100001111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001101111111011110111000101111011111111111111010001100101011000111,
	240'b101010011100101011111111111011011011010110101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111010110110101111101010001011110011110101111111111011011110111100,
	240'b101011111101011011111111110010011010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001110001011110111111110100110011111010011011010110111111111100001011000101,
	240'b101111101110001111111111101111101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011110111101101111011010101111110001011101111001001111111111101001111001011,
	240'b101111111110010011111111101111101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101011111111000001111100001100110111001000111111111101010111001100,
	240'b101111111110010011111111101111101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001110101001111100111111001111111101100110111001000111111111101010111001100,
	240'b101111111110010011111111101111101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110111111101111100110111000010111110011100111011001000111111111101010111001100,
	240'b101111111110010011111111101111101010100010101010101010011010100010101000101010001010100110101001101010101010101010101010101010101010101010101010101010101010100011000000111101111010111110100110111011001100111011001000111111111101010111001100,
	240'b101111111110010011111111101111101010011110101000101100111011111111000000101111011011010010101101101010001010100010101001101010101010101010101010101010101010100110110100111101011101101011010000111110011011111011001001111111111101010111001100,
	240'b101111111110010011111111101111101010100111010000111101001111110011111100111110111111011111101011110110001100000110101110101010001010100110101010101010101010101010101001110010101111011011111000110101101010100011001011111111111101010111001101,
	240'b101111111110010011111111101111011101001011111111111111111111111111111111111111111111111111111111111111111111110111101011110010101010111010101000101010101010101010101010101010011011001110110110101010101010011011001011111111111101010111001101,
	240'b101111111110010011111111110100011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110111110101010001010100110101010101010101010100110101001101010101010011111001011111111111101010111001101,
	240'b101111111110010011111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111010101010101001101010101010101010101010101010101010011111001011111111111101010111001101,
	240'b101111111110001111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111011111111111111111111111101101100010101011101010011010101010101010101010101010011111001011111111111101010111001100,
	240'b101111111110001111111111111110111111111111111111111111111111111111111111111111111111111111111111111100101101000011000000110000101101011011110111111111111111111111011001101010111010100110101010101010101010011111001011111111111101010111001100,
	240'b101111111110001111111111111110001111111111111111111111111111111111111111111111111111111111101010101101011010011110100110101001101010011110111100111100111111111111111111110100101010100010101010101010101010011111001011111111111101010111001100,
	240'b101111111110001111111111111101001111111111111111111111111111111111111111111111111111100010110111101001101010101010110101101101001010100110100110110001001111110111111111111110111100001010101000101010101010011111001011111111111101010111001100,
	240'b101111111110010011111111111010111111111111111111111111111111111111111111111111111111100011001100101011111101001111110111111101101100110010101000101010111110100111111111111111111111000010110001101010011010011111001011111111111101010111001100,
	240'b101111111110010011111110111000011111111111111111111111111111111111111111111111111111111111111111111011111111111011111111111111111111100110110101101001101101011011111111111111111111111111010110101010001010011111001011111111111101010111001100,
	240'b101111111110010011111111110100101111101111111111111111111111111111111111111111111111111111111111111111111110111011011110110111111111000011000001101001011100111011111111111111111111111111111000101101111010010111001011111111111101010111001101,
	240'b101111111110010011111111110001101111000111111111111111111111111111111111111111111111111111111001110011011010111010101000101010001011000110110000101001111100110111111111111111111111111111111111110110001010010111001011111111111101010111001101,
	240'b101111111110010011111111101111011101111011111111111111111111111111111111111111111111111011001100101001111010011110101000101010001010100010101001101001111100110111111111111111111111111111111111111101001010111111001010111111111101010111001101,
	240'b101111111110010011111111101111001100010111111111111111111111111111111111111111111110100110101100101010001011110111011111110111001011011110101001101001111100110111111111111111111111111111111111111111111100010011001000111111111101010111001101,
	240'b101111111110010011111111101111011010111011110010111111111111111111111111111111111101000010100101101101011111010011111111111111111110101110101110101001111100110111111111111111111111111111111111111111111101110011001010111111111101010111001101,
	240'b101111111110010011111111101111101010010111010100111111111111111111111111111111111100010010100101110010101111111111111111111111111111111010111110101001011100110111111111111111111111111111111111111111111110111011010000111111111101010111001100,
	240'b101111111110010011111111101111101010011010110011111101001111111111111111111111111100010010100101110010101111111111111111111111111111110110111110101001011101000011111111111111111111111111111111111111111111100011011011111111111101010111001100,
	240'b101111111110010011111111101111101010100010101000110011101111111111111111111111111101000010100110101101001111001111111111111111111110100110101110101001111101110111111111111111111111111111111111111111111111110111100110111111111101010111001100,
	240'b101111111110010011111111101111101010100010101001101011001110011111111111111111111110101010101100101010001011101111011110110110101011011010100111101100101111010011111111111111111111111111111111111111111111111011110001111111111101010111001100,
	240'b101111111110010011111111101111101010100010101010101010001011100011110101111111111111111011001111101001111010011110101000101010001010011110101001110110101111111111111111111111111111111111111111111111111111111111111000111111111101010111001100,
	240'b101111111110010011111111101111101010100010101010101010101010100011000100111110101111111111111011110100011011000110101010101010101011010011011001111111101111111111111111111111111111111111111111111111111111111111111100111111111101010111001100,
	240'b101111111110010011111111101111101010100010101010101010101010101010101000110010011111101111111111111110011110000011010001110100111110010011111011111111111111111111111111111111111111111111111111111111111111111111111110111111111101010111001101,
	240'b101111111110010011111111101111101010100010101010101010101010101010101010101010001100011011111000111001001011101010111101101111001011110011101011111111111111111111111111111111111111111111111111111111111111111111110110111111111101010111001101,
	240'b101111111110010011111111101111101010100010101010101010101010101010101010101010101010100010111100111001001111010111110101111101001111010011111100111111111111111111111111111111111111111111111111111111111111101111100001111111111101010111001101,
	240'b101111111110010011111111101111101010100010101000101010001010100010101001101010101010101010101000101011111101000111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111001100111111111101010111001101,
	240'b101111111110010011111111101111101010011110111011110101111100101110101101101010011010101010101010101010011010100010110100110100001110110111111100111111111111111111111111111111111111111111111111111010101011001011001001111111111101010111001101,
	240'b101111111110010011111111101111011011011111110101111100101111101011010111101010011010101010101010101010101010101010101001101010001010111110111101110011101101110111100101111010011110011011010001101100011010010111001011111111111101010111001100,
	240'b101111111110010011111111101111001101011011101011101011111100101011110101101100101010100110101010101010101010101010101010101010101010100110101000101010001010100010101010101011001010101010101000101010011010011111001011111111111101010111001100,
	240'b101111111110010011111111101111001101111011100011101001011011111111110110101101011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010011111001011111111111101010111001100,
	240'b101111111110010011111111101111001101110011111101110111111111000111100101101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111001011111111111101010111001100,
	240'b101111111110010011111111101111001101110111110011111010101110000010110100101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111001011111111111101010111001100,
	240'b101111111110010011111111101111001101011011101011101100101011111110111011101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111001011111111111101010111001100,
	240'b101110011101111011111111101111111011011111110110111100101111101011010100101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111001101111111111100111011001001,
	240'b101001111100111111111111110101111010011010111010110101011100100110101100101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010101011100011111111111011100111000000,
	240'b101100101100001111111111111110101100111110111000101101111011011110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110101101011111111101111110101011101110111010,
	240'b111010101101000011011010111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111110100001101110011011100,
	240'b111111101111011110111101110101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011001110110010101111110111111011,
	240'b111100011111010111111001110000001010000010101000101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101011101010111010101110101011101001111001111011000001111100101111000111110011,
	240'b111101111111100011101101101100111010010010111001101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101101101010001110111111111100101111011111110111,
	240'b111111111111111111011001101101101011110111010101110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110100101011101111000000111011111111111111111101,
	240'b111111101110100010111101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101111111111010011110100,
	240'b110100011100010111110010111111111101101010100101101000001010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011010000110100001101000011001111010011101101010011110010111111111111010001100101011000111,
	240'b101010011100101011111111110010010010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010000000000000011010111100000111111111011011110111100,
	240'b101011111101011111111111010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001101000011011110011011100000000010000100111111111100001011000101,
	240'b101111101110001111111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100110111001101110000001111010110011001101011101111111111101010011001011,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010100000001000011110100010110101001011001111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111101110111011101100111110110110101001011001111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000111010000110101001001001111011000110110101011001111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001111001100000111100000000110001100110111001011001111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000110100011111101000010001110000001110100001000000000000000000000000000000000000000000000000000000000000000000000011110111000101001000001110001111011000011101001011100111111111101010111001100,
	240'b101111111110010011111111001110110000001101110010110111011111011011110111111100101110011011000011100010100100010100001011000000000000000000000000000000000000000000000000010111111110001111101011100001010000000101100010111111111101010111001101,
	240'b101111111110010011111111001110100111100111111111111111111111111111111111111111111111111111111111111111111111100111000100011000100000110000000000000000000000000000000000000000000001110000100100000000000000000001100011111111111101010111001101,
	240'b101111111110010011111010011101001110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110100111011000000000000000000000000000000000000000000000000000000000000000001100011111111111101010111001101,
	240'b101111111110010011111010110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011011110000001100000000000000000000000000000000000000000000000001100011111111111101010111001101,
	240'b101111111110010011111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110101111111111111111111111011000100100000110000000000000000000000000000000000000000001100011111111111101010111001100,
	240'b101111111110001111111111111101001111111111111111111111111111111111111111111111111111111111111111110110010111001101000010010001111000001111100111111111111111111110001110000001010000000000000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111111111011001111111111111111111111111111111111111111111111111111111111000001001000110000000000000000000000000000000000111000110110101111111111111110011101110000000000000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111101110111101111111111111111111111111111111111111111111111111110101000101001000000000000000000100010000111100000000000000000010011101111100011111111111100110100100000000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111001110000111111111111111111111111111111111111111111111111111110101101100110000100010111110011101000111000110110011000000000000001011011111011111111111111111101001000010111000000000000000001100011111111111101010111001100,
	240'b101111111110010011110111101001001111111011111111111111111111111111111111111111111111111111111110110011111111110011111111111111111110110100100010000000001000001111111111111111111111111110000101000000000000000001100011111111111101010111001100,
	240'b101111111110010011111010011110001111001011111111111111111111111111111111111111111111111111111111111111111100110110011100101000001101000101000101000000000110101111111111111111111111111111101001001010000000000001100011111111111101010111001101,
	240'b101111111110010011111101010100101101011011111111111111111111111111111111111111111111111111101110011010000000111100000000000000000001010100010010000000000110100011111111111111111111111111111111100010010000000001100011111111111101010111001101,
	240'b101111111110010011111111001110101001110011111111111111111111111111111111111111111111101101100110000000000000000000000000000000000000000000000000000000000110100011111111111111111111111111111111110111010000111101011111111111111101010111001101,
	240'b101111111110010011111111001101100101000111111110111111111111111111111111111111111011111000000110000000000011101010011111100101010010100000000000000000000110100011111111111111111111111111111111111111100100110101011011111111111101010111001101,
	240'b101111111110010011111111001110100000110111011000111111111111111111111111111111110111000100000000001000011101111011111111111111111100001000001110000000000110100011111111111111111111111111111111111111111001011001011111111111111101010111001101,
	240'b101111111110010011111111001111010000000001111110111111111111111111111111111111100100110100000000011000001111111111111111111111111111101100111101000000000110100011111111111111111111111111111111111111111100110001110010111111111101010111001100,
	240'b101111111110010011111111001111100000000000011011110111101111111111111111111111100100111000000000010111111111111111111111111111111111101000111100000000000111001011111111111111111111111111111111111111111110101010010011111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000011010111111111011111111111111110111001100000000000111111101101011111111111111111011111000001101000000001001101011111111111111111111111111111111111111111111100010110100111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000010011011011011111111111111111100000100001000000000000011010010011101100100010010001100000000000110011101110111111111111111111111111111111111111111111111101111010100111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000000000010101111100000111111111111110001101111000000000000000000000000000000000000000000000010100100001111111111111111111111111111111111111111111111111111110111101100111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000000000000000001001110111100001111111111110011011101000001100000000000000000010010000010001101111111001111111111111111111111111111111111111111111111111111111011110111111111111101010111001100,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000010111011111001011111111111011001010000101110110011110101010110111110101111111111111111111111111111111111111111111111111111111111111111111111011111111111101010111001101,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000101010011101010101011010011000000110111001101100011010111000011111111111111111111111111111111111111111111111111111111111111110111100011111111111101010111001101,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000000000000111000101011101101111111100001110111011101110111110101111111111111111111111111111111111111111111111111111111111111001010100101111111111101010111001101,
	240'b101111111110010011111111001111100000000000000000000000000000000000000000000000000000000000000000000100000111011011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111010010001101000111111111101010111001101,
	240'b101111111110010011111111001111100000000000110100100001110110001100001000000000000000000000000000000000000000000000100001011100101100100111110101111111111111111111111111111111111111111111111111110000010001101101011110111111111101010111001101,
	240'b101111111110010011111111001110010010100111100001110110011110111110000110000000010000000000000000000000000000000000000000000000000000111000111010011011011001100010110010101111001011010101110110000101010000000001100011111111111101010111001100,
	240'b101111111110010011111111001101101000010011000011000101000110000111100001000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000100000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111111001101111001111010101011000000000011111011100101000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111111001101111001011111111000101000001101010110110000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111111001101111001100111011011110000011010001100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011111111111101010111001100,
	240'b101111111110010011111111001101011000010111000010000110000100000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100010111111111101010111001100,
	240'b101110011101111111111111010000000010100111100011110110001111000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101010111111111100111011001001,
	240'b101001111100111111111111100010000000000000110000100000000101110000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101100111111111011100111000000,
	240'b101100101100001111111111111100010111000100101010001010000010011100101100001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101101001100111000100011111010111110101011101110111010,
	240'b111010101101000011011010111111111111111111101110111010111110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111100001111111111111111110100001101110011011100,
	240'b111111101111011110111101110101101111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111001110110010101111110111111011,
	240'b111100011111010111111001110000001010000010101000101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101011101010111010101110101011101001111001111011000001111100101111000111110011,
};
assign data = picture[addr];
endmodule