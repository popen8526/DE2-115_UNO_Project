module green_three(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100101111101011110001101100111010110110110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011010101010110001111010111111001111110101,
	240'b111011111111101111010111101111111101001111100110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001101100111010111010110011111111000011110011,
	240'b111100011101001111001101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111101001011110011,
	240'b110010101100001111111101111111111101010010110011101100011011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011000010101110101101001101101011111111111110011011111011001000,
	240'b100110001110000111111111110000000101101001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110101101101100111010100000101111111001110111111111101001010100011,
	240'b101010001110111111111010011110100100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011010111101100111110101101010010100111010001000111111111110011110110101,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000101001001110010010100101110011110101111001111000111110111110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100110111110101010011001011001100101001001111010111110111110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101010011111110111011100010111100100111001111010111110111110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010011010000101011101010101000101000001111010111110111110111010111011,
	240'b101110001110111111110010011011010101001001010100010100010100111101001111010100000101001001010011010101000101010101010101010101010101010101010101010101010101001001110000111011110111011101001001101001001001110001110111111110111110111010111011,
	240'b101110001110111111110010011011010100111101010110011101111000111110001110100001100111010101100001010101010101000001010011010101010101010101010101010101010101010001011101110110011101001010100111111101101001011001110101111110111110111010111011,
	240'b101110001110111111110010011010100110000110111110111101011111111111111111111111001111001111100101110000101001010001100101010100010101001001010101010101010101010101010010011110101101100111101111101100010101011001111001111110111110111010111011,
	240'b101110001110111111110001011101001100100011111111111111111111111111111111111111111111111111111111111111111111111111100110101011010110100101010001010101000101010101010101010100100101101101100010010101010101000001111010111110111110111010111011,
	240'b101110001110111111101101101011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010010100010101010101001101010101010101010101010001010011010101000101000101111010111110111110111010111011,
	240'b101110001110111011110001111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101110101111001010010010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111011111000111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111101001111111111111111111111111100110101100100010100010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110110111111001111100111111111111111111111111111111111111111111111111111111111111111111111011111001111001110001011100111010011111110101111111111111111111010000011000110101001001010101010101010101000101111010111110111110111010111011,
	240'b101110001110111011110111111100001111111111111111111111111111111111111111111111111111111111110111100010000100111001001110010011100100111110010111111110111111111111111111110001010101101001010011010101010101000101111010111110111110111010111011,
	240'b101110001110111011110100111010111111111111111111111111111111111111111111111111111111111111000110010100110101010001110011011011110101000101010110110101001111111111111111111111111010011101010001010101010101000101111010111110111110111010111011,
	240'b101110001110111011101111110111101111111111111111111111111111111111111111111111111111111110011111010010110111000011101110111000110111000001011100101110001111111111111111111111111111010101111101010100010101000101111010111110111110111010111011,
	240'b101110001110111111101110110001101111111111111111111111111111111111111111111111111111111110011100010010110111010111111001111111111110100111100001111100001111111111111111111111111111111111010001010110010100111101111010111110111110111010111011,
	240'b101110001110111111101101101001011111110111111111111111111111111111111111111111111111111110111111010100110101011010000101100111001101110011111111111111111111111111111111111111111111111111111101100011110100110001111010111110111110111010111011,
	240'b101110001110111111101111100001101110111111111111111111111111111111111111111111111111111111011100010111100101001101010000010011011011110011111111111111111111111111111111111111111111111111111111110101000101010101111001111110111110111010111011,
	240'b101110001110111111110001011011111100110111111111111111111111111111111111111111111111011110000111010100100101000101011001010111101100001011111111111111111111111111111111111111111111111111111111111110100111101101110110111110111110111010111011,
	240'b101110001110111111110010011001111001100111111111111111111111111111111111111111111100010001010011010100101000110011010010110111011111001011111111111111111111111111111111111111111111111111111111111111111010111101110110111110111110111010111011,
	240'b101110001110111111110010011010100110010111101100111111111111111111111111111111111001000101001100011100111111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010000011111110011110111010111011,
	240'b101110001110111111110010011011010100111010110000111111111111111111111111111111000111111101001011100110101111111111111111111111111111111111100100110100111110001111111111111111111111111111111111111111111111001110011100111101111110111010111011,
	240'b101110001110111111110010011011010100111101101011111011001111111111111111111111101000001101001011100100011111111111111111111111111111111010000101010100101001011111111111111111111111111111111111111111111111111010111010111101101110111010111011,
	240'b101110001110111111110010011011010101001001010001100111111111111111111111111111111010000001001101011000111101100111111111111111111100110001011011010011011011001011111111111111111111111111111111111111111111111111010100111101111110111010111011,
	240'b101110001110111111110010011011010101001001010011010110101100111111111111111111111101100101011100010100000110100110100011100111110110001101001111011001001110011011111111111111111111111111111111111111111111111111101010111110001110111010111011,
	240'b101110001110111111110010011011010101001001010101010100010110111111100111111111111111111010101001010100100100111101001111010011110100111101010110101110001111111111111111111111111111111111111111111111111111111111110011111110011110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101000010000010111100001111111111111011101100110110110101011011010111000111001010111111111111101111111111111111111111111111111111111111111111111111111111110101111110101110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010000100001111110111011111111111111111111000011010111110110011111001111111111111111111111111111111111111111111111111111111111111111111111111111110101111110101110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010100000111110111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111110001110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101000101101010101111101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111010111101101110111010111011,
	240'b101110001110111111110010011011010101000101010001010100100101000101010100010101010101010101010010010101011000100111010010111111011111111111111111111111111111111111111111111111111111111111111111111111111100111110000011111110011110111010111011,
	240'b101110001110111111110010011011000101001110011000110011101010101101011111010101000101010101010101010101000101000001011011100010001100001111101000111111011111111111111111111111111111111111111111110101100110101101110110111110111110111010111011,
	240'b101110001110111111110010011010011001001011110110110011111111000010110101010100110101010101010101010101010101010101010100010100000101010001100111100000011001110010110000101110101011011110010010010111110100111001111010111110111110111010111011,
	240'b101110001110111111110001011011011011110010110100010011001001010111100111011000110101001101010101010101010101010101010101010101010101010001010011010100010101000001010000010100000101000001010000010100110101000101111010111110111110111010111011,
	240'b101110001110111111110010011011010101110101011001010011101001100111100110011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111111110010011011010100111001101000110010011111000110101110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111111110010011011010101000001101000110001101111011110000011010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111111110010011010100110011010111000100000001110100010010111010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111001111110111110111010111011,
	240'b101011101111000011110111011100010101101011010100111110101110011001101111010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110000001111111101110101010111000,
	240'b100101101110011111111111101010000100111001100001100010110110110101001110010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110101001110111000111111111101011110100101,
	240'b101101111100101011111111111110001011000010001001100001111000100110001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001011100111111011111111111100001010110110,
	240'b111011001100011011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111100011011101101,
	240'b111110001111001111000000110011101110110011111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110100111001100110001101111010111111000,
	240'b111111111111011011101010101010011001100010101111101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101011011001100010111011111111011111111111111011,
	240'b111100101111101011110001101100111010110110110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011010101010110001111010111111001111110101,
	240'b111011111111101111010111101111111101001111100110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001011100111010111010110011111111000011110011,
	240'b111100011101001111001101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111101001011110011,
	240'b110010101100001111111101111111111110100111011001110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101011111010111110110011110110111111111111110011011111011001000,
	240'b100110001110000111111111110111111010110110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111010110110110011101010001010111111100111111111111101001010100011,
	240'b101010001110111011111101101111001010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101101011110110011111010110101001010011011000100111111111110011010110101,
	240'b101110001110111011111010101101101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110100101111000111010010111001111010111110111011111111101110111010111011,
	240'b101110001110111011111010101101101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110011011111010011001100101100101010100110111100111111101110111010111011,
	240'b101110001110111011111010101101101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110101001111111011101110101011111010011110111100111111101110111010111011,
	240'b101110001110111011111010101101101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110011111101001101000010101110101010101010100010111100111111101110111010111011,
	240'b101110001110111011111010101101101010100110101010101010001010011110100111101010001010100010101001101010101010101010101010101010101010101010101010101010101010100010111000111101111011101110100100110100101100111010111011111111101110111010111011,
	240'b101110001110111011111010101101101010011110101010101110111100011111000111110000101011101010110000101010101010011110101001101010101010101010101010101010101010100110101110111011001110100111010011111110111100101110111010111111101110111010111011,
	240'b101110001110111011111010101101001011000011011111111110101111111111111111111111011111100111110010111000001100100110110010101010001010100110101010101010101010101010101000101111001110110011110111110110001010101110111100111111101110111010111011,
	240'b101110001110111011111001101110011110010011111111111111111111111111111111111111111111111111111111111111111111111111110011110101101011010010101000101010101010101010101010101010011010110110110001101010101010011110111100111111101110111010111011,
	240'b101110001110111011110111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011001001101010101010100110101010101010101010100110101001101010101010100010111100111111101110111010111011,
	240'b101110001110110111111001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111010111110101001101010101010101010101010101010101010100010111100111111101110111010111011,
	240'b101110001110110111111100111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111110101111111111111111111111111110011010110010101010001010101010101010101010101010100010111100111111101110111010111011,
	240'b101110001110110111111101111110011111111111111111111111111111111111111111111111111111111111111111111101111100111010111000101110011101001111111010111111111111111111100111101100011010100110101010101010101010100010111100111111101110111010111011,
	240'b101110001110110111111100111101111111111111111111111111111111111111111111111111111111111111111011110001001010011010100111101001111010011111001011111111011111111111111111111000101010110010101001101010101010100010111100111111101110111010111011,
	240'b101110001110110111111010111101011111111111111111111111111111111111111111111111111111111111100010101010011010100110111001101101111010100010101010111010101111111111111111111111111101001110101000101010101010100010111100111111101110111010111011,
	240'b101110001110111011111000111011111111111111111111111111111111111111111111111111111111111111001111101001011011011111110111111100011011100010101101110111001111111111111111111111111111101010111110101010001010100010111100111111101110111010111011,
	240'b101110001110111011110111111000101111111111111111111111111111111111111111111111111111111111001110101001011011101011111100111111111111010011110000111110001111111111111111111111111111111111101000101011001010011110111100111111101110111010111011,
	240'b101110001110111011110111110100011111111011111111111111111111111111111111111111111111111111011111101010011010101011000010110011011110110111111111111111111111111111111111111111111111111111111110110001111010010110111100111111101110111010111011,
	240'b101110001110111011111000110000101111011111111111111111111111111111111111111111111111111111101110101011111010100110100111101001101101110111111111111111111111111111111111111111111111111111111111111010011010101010111100111111101110111010111011,
	240'b101110001110111011111001101101111110011011111111111111111111111111111111111111111111101111000011101010001010100010101100101011101110000011111111111111111111111111111111111111111111111111111111111111011011110110111010111111101110111010111011,
	240'b101110001110111011111001101100111100110011111111111111111111111111111111111111111110000110101001101010011100010111101000111011101111100011111111111111111111111111111111111111111111111111111111111111111101011110111010111111101110111010111011,
	240'b101110001110111011111010101101001011001011110110111111111111111111111111111111111100100010100101101110011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111000001111111011110111010111011,
	240'b101110001110111011111010101101101010011111011000111111111111111111111111111111011011111110100101110011001111111111111111111111111111111111110001111010011111000111111111111111111111111111111111111111111111100111001101111111001110111010111011,
	240'b101110001110111011111010101101101010011110110101111101011111111111111111111111101100000110100101110010001111111111111111111111111111111011000010101010001100101111111111111111111111111111111111111111111111111011011100111110111110111010111011,
	240'b101110001110111011111010101101101010100010101000110011111111111111111111111111111101000010100110101100011110110011111111111111111110010110101101101001101101100011111111111111111111111111111111111111111111111111101010111111001110110110111011,
	240'b101110001110111011111010101101101010100110101001101011001110011111111111111111111110110010101101101010001011010011010001110011111011000110100111101100011111001011111111111111111111111111111111111111111111111111110100111111001110110110111011,
	240'b101110001110111011111010101101101010100110101010101010001011011111110011111111111111111111010100101010001010011110100111101001111010011110101011110111001111111111111111111111111111111111111111111111111111111111111001111111011110110110111011,
	240'b101110001110111011111010101101101010100110101010101010101010100011000000111101111111111111111101110110011011011010101101101011101011100011011111111111111111111111111111111111111111111111111111111111111111111111111010111111011110110110111011,
	240'b101110001110111011111010101101101010100110101010101010101010101010101000110000111111011111111111111111111111011111101011111011001111100111111111111111111111111111111111111111111111111111111111111111111111111111111010111111101110110110111011,
	240'b101110001110111011111010101101101010100110101010101010101010101010101010101010001011111011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111111001110110110111011,
	240'b101110001110111011111010101101101010100110101010101010101010101010101010101010101010100010110100110111101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011101111110111110111010111011,
	240'b101110001110111011111010101101101010100110101000101010011010100010101001101010101010101010101000101010101100010011101001111111101111111111111111111111111111111111111111111111111111111111111111111111111110011111000001111111011110111010111011,
	240'b101110001110111011111010101101101010100111001011111001111101010110101111101010011010101010101010101010101010100010101101110001001110000111110011111111101111111111111111111111111111111111111111111010101011010110111011111111101110111010111011,
	240'b101110001110111011111001101101001100100111111011111001111111100011011010101010011010101010101010101010101010101010101001101010001010100110110011110000001100110111011000110111011101101111001001101011111010011010111100111111101110111010111011,
	240'b101110001110111011111001101101101101111011011001101001101100101011110011101100011010100110101010101010101010101010101010101010101010101010101001101010001010100010101000101010001010100010101000101010011010100010111100111111101110111010111011,
	240'b101110001110111011111010101101101010111010101100101001101100110011110010101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111100111111101110111010111011,
	240'b101110001110111011111010101101101010011110110100111001001111100011010110101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111100111111101110111010111011,
	240'b101110001110111011111010101101101010100010110100111000101111101111000001101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111100111111101110111010111011,
	240'b101110001110111011111010101101001011001111011100101111111111010011001011101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111100111111101110111010111011,
	240'b101011101110111111111100101110001010110011101010111111001111001010110111101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011111000000111111111110101010111000,
	240'b100101101110011011111111110100111010011010110000110001011011011010100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010100111011100111111111101011110100101,
	240'b101101111100101011111111111110111101011111000100110000111100010011000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001101101110011111101111111111100001010110110,
	240'b111011001100011011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111100011011101101,
	240'b111110001111001111000000110011101110110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110111110100111001100110001101111010111111000,
	240'b111111111111011011101010101010011001100010101111101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101011011001100010111011111111011111111111111011,
	240'b111100101111101011110001101100111010110110110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011010101010110001111010111111001111110101,
	240'b111011111111101111010111101111111101001111100110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001101100111010111010110011111111000011110011,
	240'b111100011101001111001101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111101001011110011,
	240'b110010101100001111111101111111111101010010110011101100011011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011000010101110101101001101101011111111111110011011111011001000,
	240'b100110001110000111111111110000000101101001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010011110101101101100111010100000101111111001110111111111101001010100011,
	240'b101010001110111111111010011110100100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011010111101100111110101101010010100111010001000111111111110011110110101,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000101001001110010010100101110011110101111001111000111110111110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100110111110101010011001011001100101001001111010111110111110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101010011111110111011100010111100100111001111010111110111110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010011010000101011101010101000101000001111010111110111110111010111011,
	240'b101110001110111111110010011011010101001001010100010100010100111101001111010100000101001001010011010101000101010101010101010101010101010101010101010101010101001001110000111011110111011101001001101001001001110001110111111110111110111010111011,
	240'b101110001110111111110010011011010100111101010110011101111000111110001110100001100111010101100001010101010101000001010011010101010101010101010101010101010101010001011101110110011101001010100111111101101001011001110101111110111110111010111011,
	240'b101110001110111111110010011010100110000110111110111101011111111111111111111111001111001111100101110000101001010001100101010100010101001001010101010101010101010101010010011110101101100111101111101100010101011001111001111110111110111010111011,
	240'b101110001110111111110001011101001100100011111111111111111111111111111111111111111111111111111111111111111111111111100110101011010110100101010001010101000101010101010101010100100101101101100010010101010101000001111010111110111110111010111011,
	240'b101110001110111111101101101011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010010100010101010101001101010101010101010101010001010011010101000101000101111010111110111110111010111011,
	240'b101110001110111011110001111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101110101111001010010010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111011111000111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111101001111111111111111111111111100110101100100010100010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110110111111001111100111111111111111111111111111111111111111111111111111111111111111111111011111001111001110001011100111010011111110101111111111111111111010000011000110101001001010101010101010101000101111010111110111110111010111011,
	240'b101110001110111011110111111100001111111111111111111111111111111111111111111111111111111111110111100010000100111001001110010011100100111110010111111110111111111111111111110001010101101001010011010101010101000101111010111110111110111010111011,
	240'b101110001110111011110100111010111111111111111111111111111111111111111111111111111111111111000110010100110101010001110011011011110101000101010110110101001111111111111111111111111010011101010001010101010101000101111010111110111110111010111011,
	240'b101110001110111011101111110111101111111111111111111111111111111111111111111111111111111110011111010010110111000011101110111000110111000001011100101110001111111111111111111111111111010101111101010100010101000101111010111110111110111010111011,
	240'b101110001110111111101110110001101111111111111111111111111111111111111111111111111111111110011100010010110111010111111001111111111110100111100001111100001111111111111111111111111111111111010001010110010100111101111010111110111110111010111011,
	240'b101110001110111111101101101001011111110111111111111111111111111111111111111111111111111110111111010100110101011010000101100111001101110011111111111111111111111111111111111111111111111111111101100011110100110001111010111110111110111010111011,
	240'b101110001110111111101111100001101110111111111111111111111111111111111111111111111111111111011100010111100101001101010000010011011011110011111111111111111111111111111111111111111111111111111111110101000101010101111001111110111110111010111011,
	240'b101110001110111111110001011011111100110111111111111111111111111111111111111111111111011110000111010100100101000101011001010111101100001011111111111111111111111111111111111111111111111111111111111110100111101101110110111110111110111010111011,
	240'b101110001110111111110010011001111001100111111111111111111111111111111111111111111100010001010011010100101000110011010010110111011111001011111111111111111111111111111111111111111111111111111111111111111010111101110110111110111110111010111011,
	240'b101110001110111111110010011010100110010111101100111111111111111111111111111111111001000101001100011100111111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010000011111110011110111010111011,
	240'b101110001110111111110010011011010100111010110000111111111111111111111111111111000111111101001011100110101111111111111111111111111111111111100100110100111110001111111111111111111111111111111111111111111111001110011100111101111110111010111011,
	240'b101110001110111111110010011011010100111101101011111011001111111111111111111111101000001101001011100100011111111111111111111111111111111010000101010100101001011111111111111111111111111111111111111111111111111010111010111101101110111010111011,
	240'b101110001110111111110010011011010101001001010001100111111111111111111111111111111010000001001101011000111101100111111111111111111100110001011011010011011011001011111111111111111111111111111111111111111111111111010100111101111110111010111011,
	240'b101110001110111111110010011011010101001001010011010110101100111111111111111111111101100101011100010100000110100110100011100111110110001101001111011001001110011011111111111111111111111111111111111111111111111111101010111110001110111010111011,
	240'b101110001110111111110010011011010101001001010101010100010110111111100111111111111111111010101001010100100100111101001111010011110100111101010110101110001111111111111111111111111111111111111111111111111111111111110011111110011110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101000010000010111100001111111111111011101100110110110101011011010111000111001010111111111111101111111111111111111111111111111111111111111111111111111111110101111110101110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010000100001111110111011111111111111111111000011010111110110011111001111111111111111111111111111111111111111111111111111111111111111111111111111110101111110101110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010100000111110111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111110001110111010111011,
	240'b101110001110111111110010011011010101001001010101010101010101010101010101010101010101000101101010101111101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111010111101101110111010111011,
	240'b101110001110111111110010011011010101000101010001010100100101000101010100010101010101010101010010010101011000100111010010111111011111111111111111111111111111111111111111111111111111111111111111111111111100111110000011111110011110111010111011,
	240'b101110001110111111110010011011000101001110011000110011101010101101011111010101000101010101010101010101000101000001011011100010001100001111101000111111011111111111111111111111111111111111111111110101100110101101110110111110111110111010111011,
	240'b101110001110111111110010011010011001001011110110110011111111000010110101010100110101010101010101010101010101010101010100010100000101010001100111100000011001110010110000101110101011011110010010010111110100111001111010111110111110111010111011,
	240'b101110001110111111110001011011011011110010110100010011001001010111100111011000110101001101010101010101010101010101010101010101010101010001010011010100010101000001010000010100000101000001010000010100110101000101111010111110111110111010111011,
	240'b101110001110111111110010011011010101110101011001010011101001100111100110011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111111110010011011010100111001101000110010011111000110101110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111111110010011011010101000001101000110001101111011110000011010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111010111110111110111010111011,
	240'b101110001110111111110010011010100110011010111000100000001110100010010111010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111001111110111110111010111011,
	240'b101011101111000011110111011100010101101011010100111110101110011001101111010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110000001111111101110101010111000,
	240'b100101101110011111111111101010000100111001100001100010110110110101001110010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011110101001110111000111111111101011110100101,
	240'b101101111100101011111111111110001011000010001001100001111000100110001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001011100111111011111111111100001010110110,
	240'b111011001100011011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111100011011101101,
	240'b111110001111001111000000110011101110110011111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110111110100111001100110001101111010111111000,
	240'b111111111111011011101010101010011001100010101111101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101011011001100010111011111111011111111111111011,
};
assign data = picture[addr];
endmodule