module green_skip(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100001111001111110101101100011001110010101001101010111010101010101010101010101010101010101010101010111010101110101011101010111010101110101010101010101010101010101010101010111010101110101011101010101001111010100010111001001111001111110000,
	240'b111100001110101111000100110011101110101011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110110111010000101110101110011011110001,
	240'b111011111100000011011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001101011101011101101,
	240'b101111001100101111111111111110001011010110010010100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010000100011011000110010001110100100011010110111110010111111111101001110111101,
	240'b100111001110100011111111101010000101000001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100110101010110011110011000010101101010010011010100110110010110111111011111011010011000,
	240'b101100001111100111110110011011100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110011111001011111101011111011011110001101000010101001001100011111010011111111110101101,
	240'b101101101111110111101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101101100010111111111101010100110100110100111111101111000100101011011111000001111111010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011101101110110111011000111001000110111101001100101111111100110101011111111000001111111010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100100001110000101101100110011111110001001100100100011111101111101101010110111111111111010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001101110101101100101011000101101110111010000101100001101100001100101110111111111111010111000,
	240'b101101101111110111101110011010010101001001010011010100000100111101001111010100000101000001010001010100110101010101010101010101010101010101010011011000111110011110110010010100100110101011100110111111111010110001011011111000001111111010111000,
	240'b101101101111110111101110011010010100111101100000100100001010111010101101101000111000111101110110011000000101001001010001010101000101010101010101010100011001001011110110110100101011101011101110110110110110010001011101111000011111111010111000,
	240'b101101101111110111101110011001010111001011010111111111111111111111111111111111111111111111111000110111101011011010000000010110100101000101010100010101010101001110000100110010001101100110110000011010000101000001011111111000011111111010111000,
	240'b101101101111110111101011011110101101110111111111111111111111111111111111111111111111111111111111111111111111111111111001110100011000011001010101010100100101010101010001010100110101010001010010010100110101001101011111111000011111111010111000,
	240'b101101101111110111101010101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111100011001100101000101010101010101010101010001010101010101010101001101011111111000011111111010111000,
	240'b101101101111110011110001111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100111101001010001010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111101111110101111110001111111111111111111111111111111111111111111111111111111111111111111111111111000011100000110111111110111011111111111111111110111110000110010100000101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111101111110101111110001111111111111111111111111111111111111111111111111111111111100000100110100110111101100000010111110110110010010100110110011111111111110001100001010101000001010101010101010101001101011111111000011111111010111000,
	240'b101101101111101111110100111101111111111111111111111111111111111111111111111111111100001001100101010011110100111001001110010011100100111001001110010111101011010111111111111010110111010001010001010101010101001101011111111000011111111010111000,
	240'b101101101111110011110001111011111111111111111111111111111111111111111111110010010101101101010001010110010111100110011001100111000111110001010111010100000101011010111010111111111101011001011111010100110101001101011111111000011111111010111000,
	240'b101101101111110011101101110110111111111111111111111111111111111111101101011011100101000001010010011011001110011111111111111111111111100111000000011001000100111101100011111000101111111110101011010100100101001101011111111000011111111010111000,
	240'b101101101111110011101001110000011111111111111111111111111111111110110000010100000101001101010010010100111001001111111001111111111111111111111111110010010101101001001110100111001111111111110011011101010100111101011111111000011111111010111000,
	240'b101101101111110111101000101000001111110011111111111111111111100101111100010011100111101001111111010100000101001010011111111111001111111111111111111111111001000101001101011011011111000111111111110000000101001001011111111000011111111010111000,
	240'b101101101111110111101011011111111110110111111111111111111110100101100011010011111011011111101100011101010100111101010100101011011111111111111111111111111100100001010010010110011101101111111111111101010111001101011100111000011111111010111000,
	240'b101101101111110111101101011010011100100011111111111111111101111001011001010100101100111111111111110111100110101101001111010110001011101111111111111111111101110101011011010101001100101111111111111111111010110101011011111000001111111010111000,
	240'b101101101111110111101101011001001001001111111111111111111101111101011001010100101100111011111111111111111101001101100011010011110101110111001000111111111101110001011010010101001100110011111111111111111101111001101000110111111111111010111000,
	240'b101101101111110111101110011001100110000111100110111111111110101001100100010011111011000111111111111111111111111111000111010111000100111101100011110110011100011101010010010110101101110011111111111111111111100110001000110111001111111010111000,
	240'b101101101111110111101110011010010100111010100101111111111111101101111111010011000111110011111000111111111111111111111111101110100101011101001111011011110111101001001111011011111111001111111111111111111111111110101100110110111111111010111000,
	240'b101101101111110111101110011010010101000001100011111000111111111110110100010100000101001110110000111111111111111111111111111111111010111101011000010100100101001101001111101000011111111111111111111111111111111111001101110111111111111010111000,
	240'b101101101111110111101110011010010101001001010000100100001111110011110001011100110100111101011010101011001110111111111110111111111111000001111010010100010101000101100110111001011111111111111111111111111111111111100101111001001111110110111000,
	240'b101101101111110111101110011010010101001001010100010101101011111011111111110100000101111101001111010100110110111010001110100100010111010001011001010100010101100111000001111111111111111111111111111111111111111111110001111011001111110010111000,
	240'b101101101111110111101110011010010101001001010101010100100110001111011000111111111100101001101011010011110100111001001110010011100100111001001111011001001011111011111111111111111111111111111111111111111111111111110100111100011111110010111000,
	240'b101101101111110111101110011010010101001001010101010101010101000101110000111000011111111111100111101001000111011001100101011001000111001010011011111000001111111111111111111111111111111111111111111111111111111111110110111101001111110010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010000011100111101111011111111111111111111010111100110111001011111001011111111111111111111111111111111111111111111111111111111111111111111111111110110111100111111110010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010100010110101011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111010011111110110111000,
	240'b101101101111110111101110011010010101001001010101010101010101010001010100010101010101001001011100101000101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111101111111010111000,
	240'b101101101111110111101110011010010101001001010011010100100101100001010111010100010101010001010011010100010111000110111000111100011111111111111111111111111111111111111111111111111111111111111111111111111110001001110101110111101111111010111000,
	240'b101101101111110111101110011010010100111101100110101100101110000111011010100110000101011101010100010101010101000101010100011100011010011011010011111100101111110011111111111111111111111111111101110110010111011101011011111000011111111010111000,
	240'b101101101111110111101110011001110101111011010101111101011011010011000000111101111010100101010011010101010101010101010100010100100101000001011010011011001000010010011001101000111010010110001010010111110101000001011111111000011111111010111000,
	240'b101101101111110111101101011001001001110011111100111100111000000001001011100101111111000101110011010100100101010101010101010101010101010101010100010100100101000101010000010011110100111101010000010100110101001101011111111000011111111010111000,
	240'b101101101111110111101101011010001100110010111001101110111110111101110110010101101110000110011011010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111110111101101011010101101001110100101010101101100111011100101011100011101100110100010010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111110111101101011001001011011011010101010101000101111111010100111001011111000010000100010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111110111101110011001010111010011110001101111010111010010011110111111111101000001011010010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101011101111100011110110011100000100111010001011111001011111100111110101110010100110101101010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100101111010101111111010101011,
	240'b100110101110011111111111101011110101001001001011010111110111100101110011010101010100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101000010011110111111101111010010010111,
	240'b101111111100100111111111111110111100000010011101100110111001100110011010100111001001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111011011100011110111111111111101000011000000,
	240'b111100001100000111011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011101111101110,
	240'b111110011111010111000011110001111110001011110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111000111111010,
	240'b111111111111111111101010101001101001111010110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100111010000110100111111100011111111111111111,
	240'b111100001111001111110101101100011001110010101001101010111010101010101010101010101010101010101010101010111010101110101011101010111010101110101010101010101010101010101010101010111010101110101011101010101001111010100010111001001111001111110000,
	240'b111100001110101111000100110011101110101011111000111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110110111010000101110101110011011110001,
	240'b111011111100000011011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001101011101011101101,
	240'b101111001100101111111111111111001101101011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011000111110001101100010111000110110010001101011011111001111111111101001110111101,
	240'b100111001110100011111111110100111010100010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011010101010101111001100001010110101101001101010011011001011111111101111010110011000,
	240'b101100001111100011111011101101101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011001111100101111110101111101111111000110100001010100010110001111101001111110110101101,
	240'b101101101111101111110110101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111110001011111111110101001011010011010011111110111100010010101101111100001111110010111000,
	240'b101101101111101111110110101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111011011101100111100101011011110100101110111111110011010101111111100001111110010111000,
	240'b101101101111101111110110101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110001111111000010110101111001111111000110110010110001111110111110110100111011111111110010111000,
	240'b101101101111101111110110101101001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000110000101111010110110010101100011110111011101000110110001110110010110010111011111111110010111000,
	240'b101101101111101111110110101101001010100110101001101010001010011110100111101001111010100010101000101010011010101010101010101010101010101010101001101100011111001111011001101010001011010111110010111111111101011010101101111100001111110010111000,
	240'b101101101111101111110110101101001010011110101111110010001101011011010110110100011100011110111010101100001010100010101000101010011010101010101010101010001100100111111010111010001101110111110111111011011011001010101110111100001111110010111000,
	240'b101101101111101111110110101100101011100011101011111111111111111111111111111111111111111111111100111011111101101110111111101011001010100010101010101010101010100111000001111000111110110011010111101100111010100010101111111100001111110010111000,
	240'b101101101111101111110101101111001110111011111111111111111111111111111111111111111111111111111111111111111111111111111100111010001100001110101010101010011010101010101000101010011010101010101000101010011010100110101111111100001111110010111000,
	240'b101101101111101111110101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011011101101100101010100010101010101010101010101010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111111000111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101011110110101000101010101010101010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111111010111110111111111111111111111111111111111111111111111111111111111111111111111111111111100011110000111011111111011111111111111111111111011111000011101010001010101010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111111010111110111111111111111111111111111111111111111111111111111111111111110000110011011011011110110000101011111011011011001001111011001111111111111000110000101010100010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111111010111110111111111111111111111111111111111111111111111111111110000010110010101001111010011110100111101001111010011010100111101011111101101011111111111101011011101010101000101010101010100110101111111100001111110010111000,
	240'b101101101111101111111000111101111111111111111111111111111111111111111111111001001010110110101000101011001011110011001100110011011011111010101011101001111010101111011100111111111110101110101111101010011010100110101111111100001111110010111000,
	240'b101101101111101111110110111011011111111111111111111111111111111111110110101101101010100010101001101101011111001111111111111111111111110011100000101100011010011110110001111100001111111111010101101010001010100110101111111100001111110010111000,
	240'b101101101111101111110100111000001111111111111111111111111111111111010111101010001010100110101001101010011100100111111100111111111111111111111111111001001010110110100110110011011111111111111001101110101010011110101111111100001111110010111000,
	240'b101101101111101111110100110011111111111011111111111111111111110010111110101001101011110010111111101001111010100011001111111111101111111111111111111111111100100010100110101101101111100011111111111000001010100010101111111100001111110010111000,
	240'b101101101111101111110101101111111111011011111111111111111111010010110001101001111101101111110101101110101010011110101010110101101111111111111111111111111110001110101001101011001110110111111111111110101011100110101101111100001111110010111000,
	240'b101101101111101111110110101101001110010011111111111111111110111110101100101010001110011111111111111011111011010110100111101010111101110111111111111111111110111010101101101010101110010111111111111111111101011010101101111100001111110010111000,
	240'b101101101111101111110110101100011100100111111111111111111110111110101100101010001110011011111111111111111110100110110001101001111010111011100011111111111110110110101101101010101110011011111111111111111110111010110011111011111111110010111000,
	240'b101101101111101111110110101100111011000011110010111111111111010010110001101001111101100011111111111111111111111111100011101011101010011110110001111011001110001110101000101011001110111011111111111111111111110011000011111011101111110010111000,
	240'b101101101111101111110110101101001010011011010010111111111111110110111111101001101011110111111100111111111111111111111111110111011010101110100111101101111011110110100111101101111111100111111111111111111111111111010101111011011111110010111000,
	240'b101101101111101111110110101101001010011110110001111100011111111111011001101010001010100111010111111111111111111111111111111111111101011110101011101010011010100110100111110100001111111111111111111111111111111111100110111011111111110010111000,
	240'b101101101111101111110110101101001010100110101000110001111111111011111000101110011010011110101101110101101111011111111111111111111111011110111101101010001010100010110011111100101111111111111111111111111111111111110010111100101111110010111000,
	240'b101101101111101111110110101101001010100110101010101010101101111011111111111010001010111110100111101010011011011111000110110010001011101010101100101010001010110011100000111111111111111111111111111111111111111111111000111101101111101110111000,
	240'b101101101111101111110110101101001010100110101010101010011011000111101100111111111110010110110101101001111010011110100111101001101010011110100111101100011101111011111111111111111111111111111111111111111111111111111010111110001111101110111000,
	240'b101101101111101111110110101101001010100110101010101010101010100010111000111100001111111111110011110100011011101010110010101100101011100111001101111100001111111111111111111111111111111111111111111111111111111111111011111110101111101110111000,
	240'b101101101111101111110110101101001010100110101010101010101010101010101000101110011110111011111111111111111111101011110011111100101111100111111111111111111111111111111111111111111111111111111111111111111111111111111010111110011111101110111000,
	240'b101101101111101111110110101101001010100110101010101010101010101010101010101010001011010011100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101001111110010111000,
	240'b101101101111101111110110101101001010100110101010101010101010100110101010101010101010100010101101110100001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111011111111110010111000,
	240'b101101101111101111110110101101001010100110101001101010011010110010101011101010001010101010101001101010001011100011011011111110001111111111111111111111111111111111111111111111111111111111111111111111111111000110111010111011111111110010111000,
	240'b101101101111101111110110101101001010011110110010110110001111000011101100110010111010101110101001101010101010100010101001101110001101001111101001111110011111110111111111111111111111111111111110111011001011101110101101111100001111110010111000,
	240'b101101101111101111110110101100111010111011101011111110101101101011011111111110111101010010101001101010101010101010101010101010001010100010101100101101101100000111001100110100011101001011000100101011111010011110101111111100001111110010111000,
	240'b101101101111101111110110101100011100111011111110111110011011111110100101110010111111100010111001101010001010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100110101111111100001111110010111000,
	240'b101101101111101111110110101100111110011011011100110111011111011110111011101010101111000011001101101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111110110101101001110100111010010101010111110011111110010101110001110110011010001101001111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111110110101100101101101111101010101010011010111111101010111100101111011111000010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111110010111000,
	240'b101101101111101111110110101100101011100111111000110111101011100111001110111111111110011110101101101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111100001111110010111000,
	240'b101011101111011111111011101101111010011011000101111100101111110011111010111001011011010110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110010111101011111110110101011,
	240'b100110101110011011111111110101111010100110100101101011111011110010111001101010101010011010100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010100011001110111111101111001110010111,
	240'b101111111100100111111111111111011101111111001110110011011100110011001100110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101101110011111011111111111101000011000000,
	240'b111100001100000111011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011101111101110,
	240'b111110011111010111000011110001111110000111110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111000111111010,
	240'b111111111111111111101010101001101001111010110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100111010000110100111111100011111111111111111,
	240'b111100001111001111110101101100011001110010101001101010111010101010101010101010101010101010101010101010111010101110101011101010111010101110101010101010101010101010101010101010111010101110101011101010101001111010100010111001001111001111110000,
	240'b111100001110101111000100110011101110101011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011110110111010000101110101110011011110001,
	240'b111011111100000011011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001101011101011101101,
	240'b101111001100101111111111111110001011010110010010100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010000100011011000110010001110100100011010110111110010111111111101001110111101,
	240'b100111001110100011111111101010000101000001001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100110101010110011110011000010101101010010011010100110110010110111111011111011010011000,
	240'b101100001111100111110110011011100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110011111001011111101011111011011110001101000010101001001100011111010011111111110101101,
	240'b101101101111110111101110011010000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101101100010111111111101010100110100110100111111101111000100101011011111000001111111010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011101101110110111011000111001000110111101001100101111111100110101011111111000001111111010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100100001110000101101100110011111110001001100100100011111101111101101010110111111111111010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001101110101101100101011000101101110111010000101100001101100001100101110111111111111010111000,
	240'b101101101111110111101110011010010101001001010011010100000100111101001111010100000101000001010001010100110101010101010101010101010101010101010011011000111110011110110010010100100110101011100110111111111010110001011011111000001111111010111000,
	240'b101101101111110111101110011010010100111101100000100100001010111010101101101000111000111101110110011000000101001001010001010101000101010101010101010100011001001011110110110100101011101011101110110110110110010001011101111000011111111010111000,
	240'b101101101111110111101110011001010111001011010111111111111111111111111111111111111111111111111000110111101011011010000000010110100101000101010100010101010101001110000100110010001101100110110000011010000101000001011111111000011111111010111000,
	240'b101101101111110111101011011110101101110111111111111111111111111111111111111111111111111111111111111111111111111111111001110100011000011001010101010100100101010101010001010100110101010001010010010100110101001101011111111000011111111010111000,
	240'b101101101111110111101010101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111100011001100101000101010101010101010101010001010101010101010101001101011111111000011111111010111000,
	240'b101101101111110011110001111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100111101001010001010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111101111110101111110001111111111111111111111111111111111111111111111111111111111111111111111111111000011100000110111111110111011111111111111111110111110000110010100000101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111101111110101111110001111111111111111111111111111111111111111111111111111111111100000100110100110111101100000010111110110110010010100110110011111111111110001100001010101000001010101010101010101001101011111111000011111111010111000,
	240'b101101101111101111110100111101111111111111111111111111111111111111111111111111111100001001100101010011110100111001001110010011100100111001001110010111101011010111111111111010110111010001010001010101010101001101011111111000011111111010111000,
	240'b101101101111110011110001111011111111111111111111111111111111111111111111110010010101101101010001010110010111100110011001100111000111110001010111010100000101011010111010111111111101011001011111010100110101001101011111111000011111111010111000,
	240'b101101101111110011101101110110111111111111111111111111111111111111101101011011100101000001010010011011001110011111111111111111111111100111000000011001000100111101100011111000101111111110101011010100100101001101011111111000011111111010111000,
	240'b101101101111110011101001110000011111111111111111111111111111111110110000010100000101001101010010010100111001001111111001111111111111111111111111110010010101101001001110100111001111111111110011011101010100111101011111111000011111111010111000,
	240'b101101101111110111101000101000001111110011111111111111111111100101111100010011100111101001111111010100000101001010011111111111001111111111111111111111111001000101001101011011011111000111111111110000000101001001011111111000011111111010111000,
	240'b101101101111110111101011011111111110110111111111111111111110100101100011010011111011011111101100011101010100111101010100101011011111111111111111111111111100100001010010010110011101101111111111111101010111001101011100111000011111111010111000,
	240'b101101101111110111101101011010011100100011111111111111111101111001011001010100101100111111111111110111100110101101001111010110001011101111111111111111111101110101011011010101001100101111111111111111111010110101011011111000001111111010111000,
	240'b101101101111110111101101011001001001001111111111111111111101111101011001010100101100111011111111111111111101001101100011010011110101110111001000111111111101110001011010010101001100110011111111111111111101111001101000110111111111111010111000,
	240'b101101101111110111101110011001100110000111100110111111111110101001100100010011111011000111111111111111111111111111000111010111000100111101100011110110011100011101010010010110101101110011111111111111111111100110001000110111001111111010111000,
	240'b101101101111110111101110011010010100111010100101111111111111101101111111010011000111110011111000111111111111111111111111101110100101011101001111011011110111101001001111011011111111001111111111111111111111111110101100110110111111111010111000,
	240'b101101101111110111101110011010010101000001100011111000111111111110110100010100000101001110110000111111111111111111111111111111111010111101011000010100100101001101001111101000011111111111111111111111111111111111001101110111111111111010111000,
	240'b101101101111110111101110011010010101001001010000100100001111110011110001011100110100111101011010101011001110111111111110111111111111000001111010010100010101000101100110111001011111111111111111111111111111111111100101111001001111110110111000,
	240'b101101101111110111101110011010010101001001010100010101101011111011111111110100000101111101001111010100110110111010001110100100010111010001011001010100010101100111000001111111111111111111111111111111111111111111110001111011001111110010111000,
	240'b101101101111110111101110011010010101001001010101010100100110001111011000111111111100101001101011010011110100111001001110010011100100111001001111011001001011111011111111111111111111111111111111111111111111111111110100111100011111110010111000,
	240'b101101101111110111101110011010010101001001010101010101010101000101110000111000011111111111100111101001000111011001100101011001000111001010011011111000001111111111111111111111111111111111111111111111111111111111110110111101001111110010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010000011100111101111011111111111111111111010111100110111001011111001011111111111111111111111111111111111111111111111111111111111111111111111111110110111100111111110010111000,
	240'b101101101111110111101110011010010101001001010101010101010101010101010101010100010110101011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111010011111110110111000,
	240'b101101101111110111101110011010010101001001010101010101010101010001010100010101010101001001011100101000101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111101111111010111000,
	240'b101101101111110111101110011010010101001001010011010100100101100001010111010100010101010001010011010100010111000110111000111100011111111111111111111111111111111111111111111111111111111111111111111111111110001001110101110111101111111010111000,
	240'b101101101111110111101110011010010100111101100110101100101110000111011010100110000101011101010100010101010101000101010100011100011010011011010011111100101111110011111111111111111111111111111101110110010111011101011011111000011111111010111000,
	240'b101101101111110111101110011001110101111011010101111101011011010011000000111101111010100101010011010101010101010101010100010100100101000001011010011011001000010010011001101000111010010110001010010111110101000001011111111000011111111010111000,
	240'b101101101111110111101101011001001001110011111100111100111000000001001011100101111111000101110011010100100101010101010101010101010101010101010100010100100101000101010000010011110100111101010000010100110101001101011111111000011111111010111000,
	240'b101101101111110111101101011010001100110010111001101110111110111101110110010101101110000110011011010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111110111101101011010101101001110100101010101101100111011100101011100011101100110100010010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111110111101101011001001011011011010101010101000101111111010100111001011111000010000100010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101101101111110111101110011001010111010011110001101111010111010010011110111111111101000001011010010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111010111000,
	240'b101011101111100011110110011100000100111010001011111001011111100111110101110010100110101101010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100101111010101111111010101011,
	240'b100110101110011111111111101011110101001001001011010111110111100101110011010101010100110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101000010011110111111101111010010010111,
	240'b101111111100100111111111111110111100000010011101100110111001100110011010100111001001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111011011100011110111111111111101000011000000,
	240'b111100001100000111011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011101111101110,
	240'b111110011111010111000011110001111110001011110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111000111111010,
	240'b111111111111111111101010101001101001111010110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100111010000110100111111100011111111111111111,
};
assign data = picture[addr];
endmodule