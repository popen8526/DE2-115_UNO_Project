module crown(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 80;
localparam Y_WIDTH = 50;
parameter [0:49][79:0] picture = {
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000001111100000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000001111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000011111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000011111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000001111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000001111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000111100000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000101100000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000111100000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000001111100000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000001111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000011111110000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000011111111000000000000000000000000000000000000,
	80'b00000001111000000001111000000000000011111111000000000000011100000000011100000000,
	80'b00000001111100000001111000000000000111111111000000000000111110000000111110000000,
	80'b00000001111100000001111100000000001111111111100000000000111110000000111110000000,
	80'b00000001111100000001111100000000001111111111100000000000111110000000111110000000,
	80'b00000000111000000000111000000000011111111111110000000000011100000000011100000000,
	80'b00000000001000000000001100000000111111111111111000000000100000000000010000000000,
	80'b00000000001100000000001100000001111111111111111100000011110000000000110000000000,
	80'b00000000000100000000001111110111111111111111111111101111110000000001100000000000,
	80'b00000000000110000000001111111111111111111111111111111111110000000011100000000000,
	80'b00000000000111000000011111111111111111111111111111111111110000000111100000000000,
	80'b00000000000011110000011111111111111111111111111111111111110000011111000000000000,
	80'b00000000000011111101111111111111111111111111111111111111111001111111000000000000,
	80'b00000000000011111111111111111111111111111111111111111111111111111111000000000000,
	80'b00000000000011111111111111111111111111111111111111111111111111111110000000000000,
	80'b00000000000001111111111111111111111111111111111111111111111111111110000000000000,
	80'b00000000000001111111111111111111111111111111111111111111111111111110000000000000,
	80'b00000000000001111111111111111111111111111111111111111111111111111110000000000000,
	80'b00000000000000111111111111111111000000000000000011111111111111111100000000000000,
	80'b00000000000000111111111100111111111111111111111111111100111111111100000000000000,
	80'b00000000000000111111011111111111111111000011111111111111111011111100000000000000,
	80'b00000000000000111111111111100000000000000000000000000111111111011100000000000000,
	80'b00000000000000111111110000000000000000000000000000000000001111110100000000000000,
	80'b00000000000000011110000000000000000000000000000000000000000001111100000000000000,
	80'b00000000000000111100000000000000000000000000000000000000000000111100000000000000,
	80'b00000000000000111000000000000000000000000000000000000000000000011100000000000000,
	80'b00000000000000110000000000000000000000000000000000000000000000001100000000000000,
	80'b00000000000000010000000000000000000000000000000000000000000000001000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
	80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		// r_data = r_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		// g_data = g_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		// b_data = b_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		r_data = {8{picture[(y_cnt - y_pin)][((x_cnt - x_pin))]}};
		g_data = {8{picture[(y_cnt - y_pin)][((x_cnt - x_pin))]}};
		b_data = {8{picture[(y_cnt - y_pin)][((x_cnt - x_pin))]}};
		// r_data = 8'b0;
		// g_data = 8'b0;
		// b_data = 8'b0;
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule