module red_five(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
    240'b111100101111100011101111110010101011101110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110011010011111100011111001111110001,
    240'b111100111110100010111110110101011110100111101001111010011110100111101001111010011110100111101010111010101110101011101010111010011110100111101001111010011110100111101001111010101110101011101010111010101110011011001000101111001110100111110000,
    240'b111000111011111011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101011111011101110,
    240'b101110011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111011000010,
    240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110010010,
    240'b101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010011110,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
    240'b101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101011,
    240'b101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110010101,
    240'b101100011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010011111,
    240'b110001111101010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100000011011000,
    240'b111011111100010011011001111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110001001100110011110010,
    240'b111101111111010011000010101011111011110111000100110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100010110001110100111111011111110110,
    240'b111100101111100111101111110010111011110010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111011011110011010100111100011111001111110010,
    240'b111100111110100010111110110101011110100111101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110011111001000101111001110100111110000,
    240'b111000111011111011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101011111011101110,
    240'b101110011110011111111111111011001010111110011011100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100110011001011110010111100110011011110111111001111111111100111011000010,
    240'b101100111111111111110010011111010100111101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001010010011100111000000001111111011111110111011110101000111111101111001010010010,
    240'b101110101111111111000101010100100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011001110010101111001111110001111101101101100101101100111011101111111010011110,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011100100111100101110011101011101110001101100011111001001111111110101111,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010100110111111110011110110010101110010001100100111001001111111110110000,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100111001111100011100111111000011100001101100011111001001111111110110000,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111001111010111101100000011000010110000001011111111001011111111110110000,
    240'b110000011111111110110110010100010101010101010011010100010101000001010000010100000101000101010011010101010101010101010101010101010101010101010101010101010101001101100110111100101000011001000110100011001011010001100000111001001111111110110000,
    240'b110000011111111110110110010100010101000101100000100000011001000010001100100000100111001101100000010100110101000001010011010101010101010101010101010101010101010001011000110011111101111010100010111011011011100101011100111001011111111110101111,
    240'b110000011111111110110110010011101000001111011001111111001111111111111111111111101111001111100000101111011000111101100011010100010101001101010101010101010101010101010010011100101101001011101011110001010110010001011100111001011111111110101111,
    240'b110000011111111110110010011110111111000111111111111111111111111111111111111111111111111111111111111111111111111111100001101000010110001101010000010101000101010101010101010100100101101101100111010101110101000101011110111001011111111110101111,
    240'b110000011111111110111011110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111010001101010101000101001101010101010101010101010001010011010101000101001101011110111001011111111110101111,
    240'b110000011111111111011010111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101110101111001010001010101010101010101010101010101010101001101011110111001011111111110101111,
    240'b110000011111111111101111111111001111111111111111111111111111111111111111111111011111010111110011111100111111001111110011111100111111001111110101111101111100011101100101010100010101010101010101010101010101001101011110111001011111111110101111,
    240'b110000011111111111110100111111001111111111111111111111111111111111111111111010010111110101101111011100010111000101110001011100010111000101110000011101001101110011010100011000110101001001010101010101010101001101011110111001011111111110110000,
    240'b110000011111111111101110111110111111111111111111111111111111111111111111111000110101110001001011010011100100111001001110010011100100111101010000010101011100111011111111110001110101101001010011010101010101001101011110111001011111111110110000,
    240'b110000011111111111100110111110011111111111111111111111111111111111111111111010101000001101110110011101110111011101110111011110000110111101010101010101111100111111111111111111111010110001010010010101000101001101011110111001011111111110110000,
    240'b110000011111111111010111111101101111111111111111111111111111111111111111111111101111101111111011111110111111101111111011111110111101001001011001010101101100111111111111111111111111100010000101010100000101001101011110111001011111111110110000,
    240'b110000011111111111001001111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101011001010101101100111111111111111111111111111111011011010111110101000101011110111001011111111110110000,
    240'b110000011111111110111001110100011111111111111111111111111111111111111111111111111111111111111111111011001100011010110110101101011001110001010111010101111100111111111111111111111111111111111111100111100100111101011110111001011111111110101111,
    240'b110000011111111110110001101011111111111111111111111111111111111111111111111111111111111010111100011010110101010101001111010011110101000001010011010110001100111111111111111111111111111111111111111000100101111101011100111001011111111110101111,
    240'b110000011111111110110001100000001111110011111111111111111111111111111111111111111011111101010111010011110101000101010011010100110101001101010010010101101100111011111111111111111111111111111111111111101001000001011001111001011111111110101111,
    240'b110000011111111110110100010111001110001011111111111111111111111111111111111011100110110101001111011000011010011011000111110001111100011111000111110010001110111111111111111111111111111111111111111111111100100101011110111001001111111110101111,
    240'b110000011111111110110110010011011010100111111111111111111111111111111111110001000101001001010101101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101110110111000101111111110101111,
    240'b110000011111111110110110010011100110110111101111111111111111111111111111101010000100110101101011111100001111111111111111111111111111110011110000111100001111101011111111111111111111111111111111111111111111111110011001111000001111111110101111,
    240'b110000011111111110110110010100010101000110101101111111111111111111111111101001100100110101101101111100011111111111111111111111111101010001101011011011101101101011111111111111111111111111111111111111111111111110111101111000001111111110110000,
    240'b110000011111111110110110010100010101001001100110111000111111111111111111110000000101000101010111110001011111111111111111111111111001100101001100010111111110011111111111111111111111111111111111111111111111111111011000111001111111111110110000,
    240'b110000011111111110110110010100010101010101010000100010111111101111111111111010100110100001001111011001111011011011001111100111110101100101001110100011001111110011111111111111111111111111111111111111111111111111101001111011111111111110110000,
    240'b110000011111111110110110010100010101010101010100010101001010111011111111111111111011011001010100010100000101001101010111010100010100111101100101110111001111111111111111111111111111111111111111111111111111111111110111111101101111111110110000,
    240'b110000011111111110110110010100010101010101010101010100110101101111000100111111111111110110101111011000100101000001001111010100110111001011010000111111111111111111111111111111111111111111111111111111111111111111111100111110011111111110110000,
    240'b110000011111111110110110010100010101010101010101010101010101001001011111110001111111111111111111111000011011100010101011110000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110101111111110101111,
    240'b110000011111111110110110010100010101010101010101010101010101010101010010010111111011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101101111111110101111,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010100100101100010100001111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110111001111111111110101111,
    240'b110000011111111110110110010100010101010001010001010100000101001001010101010101010101010001010001011101111100011011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010010011111000011111111110101111,
    240'b110000011111111110110110010100000101011110000000100100010110100101010010010101010101010101010101010100010101011110000010110000011110111011111111111111111111111111111111111111111111111111111111111111001010100001011110111001001111111110101111,
    240'b110000011111111110110101010100001010100111111000111101011110001001101111010100100101010101010101010101010101010001010001010101010110110110010010101110011101001011100000111001111110011111010000100011100101010001011101111001011111111110101111,
    240'b110000011111111110110011011010011110111010100010011100011110000010110110010100100101010101010101010101010101010101010101010101000101001001010000010100010101011101100010011001110110011101011000010100010101001001011110111001011111111110110000,
    240'b110000011111111110110100010111111000100001011000010010001011110011001011010101000101010001010101010101010101010101010101010101010101010101010101010101010101010001010011010100100101001101010100010101010101001101011110111001011111111110110000,
    240'b110000011111111110110100010111011000010110001010100110111111000010100101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001011111111110110000,
    240'b110000011111111110110001011110101111100011110100111100001100000001100000010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001011111111110110000,
    240'b110000011111111110110001011111001110111010000100011010100101010101010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001011111111110110000,
    240'b101111101111111110110011011111001111011110111110101100101011011110000011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001111111111110101011,
    240'b101101111111111111010001011101111101000111011100110111001101111010010100010011110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000100111101110101111101101111101110010101,
    240'b101100011111101111111100101010000110001101011110010111100101111001011100010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010110101111001100111111111110100010011111,
    240'b110001111101010011111111111111101110000011010110110101101101011011010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111110101011111111111111011100000011011000,
    240'b111011111100010011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110001001100110011110010,
    240'b111101111111010011000010101011111011110111000100110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100010110001110100111111011111110110,
    240'b111100101111100011101111110010101011101110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110011010011111100011111001111110001,
    240'b111100111110100010111110110101011110100111101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110011111001000101111001110100111110000,
    240'b111000111011111011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101011111011101110,
    240'b101110011110011111111111111011001010111110011011100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100110011001011110010111100110011011110111111001111111111100111011000010,
    240'b101100111111111111110010011111010100111101010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001010010011100111000000001111111011111110111011110101000111111101111001010010010,
    240'b101110101111111111000101010100100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011001110010101111001111110001111101101101100101101100111011101111111010011110,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011100100111100101110011101011101110001101100011111001001111111110101111,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010100110111111110011110110010101110010001100100111001001111111110110000,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100111001111100011100111111000011100001101100011111001001111111110110000,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000111001111010111101100000011000010110000001011111111001011111111110110000,
    240'b110000011111111110110110010100010101010101010011010100010101000001010000010100000101000101010011010101010101010101010101010101010101010101010101010101010101001101100110111100101000011001000110100011001011010001100000111001001111111110110000,
    240'b110000011111111110110110010100010101000101100000100000011001000010001100100000100111001101100000010100110101000001010011010101010101010101010101010101010101010001011000110011111101111010100010111011011011100101011100111001011111111110101111,
    240'b110000011111111110110110010011101000001111011001111111001111111111111111111111101111001111100000101111011000111101100011010100010101001101010101010101010101010101010010011100101101001011101011110001010110010001011100111001011111111110101111,
    240'b110000011111111110110010011110111111000111111111111111111111111111111111111111111111111111111111111111111111111111100001101000010110001101010000010101000101010101010101010100100101101101100111010101110101000101011110111001011111111110101111,
    240'b110000011111111110111011110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111010001101010101000101001101010101010101010101010001010011010101000101001101011110111001011111111110101111,
    240'b110000011111111111011010111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101101110101111001010001010101010101010101010101010101010101001101011110111001011111111110101111,
    240'b110000011111111111101111111111001111111111111111111111111111111111111111111111011111010111110011111100111111001111110011111100111111001111110101111101111100011101100101010100010101010101010101010101010101001101011110111001011111111110101111,
    240'b110000011111111111110100111111001111111111111111111111111111111111111111111010010111110101101111011100010111000101110001011100010111000101110000011101001101110011010100011000110101001001010101010101010101001101011110111001011111111110110000,
    240'b110000011111111111101110111110111111111111111111111111111111111111111111111000110101110001001011010011100100111001001110010011100100111101010000010101011100111011111111110001110101101001010011010101010101001101011110111001011111111110110000,
    240'b110000011111111111100110111110011111111111111111111111111111111111111111111010101000001101110110011101110111011101110111011110000110111101010101010101111100111111111111111111111010110001010010010101000101001101011110111001011111111110110000,
    240'b110000011111111111010111111101101111111111111111111111111111111111111111111111101111101111111011111110111111101111111011111110111101001001011001010101101100111111111111111111111111100010000101010100000101001101011110111001011111111110110000,
    240'b110000011111111111001001111010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101011001010101101100111111111111111111111111111111011011010111110101000101011110111001011111111110110000,
    240'b110000011111111110111001110100011111111111111111111111111111111111111111111111111111111111111111111011001100011010110110101101011001110001010111010101111100111111111111111111111111111111111111100111100100111101011110111001011111111110101111,
    240'b110000011111111110110001101011111111111111111111111111111111111111111111111111111111111010111100011010110101010101001111010011110101000001010011010110001100111111111111111111111111111111111111111000100101111101011100111001011111111110101111,
    240'b110000011111111110110001100000001111110011111111111111111111111111111111111111111011111101010111010011110101000101010011010100110101001101010010010101101100111011111111111111111111111111111111111111101001000001011001111001011111111110101111,
    240'b110000011111111110110100010111001110001011111111111111111111111111111111111011100110110101001111011000011010011011000111110001111100011111000111110010001110111111111111111111111111111111111111111111111100100101011110111001001111111110101111,
    240'b110000011111111110110110010011011010100111111111111111111111111111111111110001000101001001010101101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101110110111000101111111110101111,
    240'b110000011111111110110110010011100110110111101111111111111111111111111111101010000100110101101011111100001111111111111111111111111111110011110000111100001111101011111111111111111111111111111111111111111111111110011001111000001111111110101111,
    240'b110000011111111110110110010100010101000110101101111111111111111111111111101001100100110101101101111100011111111111111111111111111101010001101011011011101101101011111111111111111111111111111111111111111111111110111101111000001111111110110000,
    240'b110000011111111110110110010100010101001001100110111000111111111111111111110000000101000101010111110001011111111111111111111111111001100101001100010111111110011111111111111111111111111111111111111111111111111111011000111001111111111110110000,
    240'b110000011111111110110110010100010101010101010000100010111111101111111111111010100110100001001111011001111011011011001111100111110101100101001110100011001111110011111111111111111111111111111111111111111111111111101001111011111111111110110000,
    240'b110000011111111110110110010100010101010101010100010101001010111011111111111111111011011001010100010100000101001101010111010100010100111101100101110111001111111111111111111111111111111111111111111111111111111111110111111101101111111110110000,
    240'b110000011111111110110110010100010101010101010101010100110101101111000100111111111111110110101111011000100101000001001111010100110111001011010000111111111111111111111111111111111111111111111111111111111111111111111100111110011111111110110000,
    240'b110000011111111110110110010100010101010101010101010101010101001001011111110001111111111111111111111000011011100010101011110000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110101111111110101111,
    240'b110000011111111110110110010100010101010101010101010101010101010101010010010111111011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101101111111110101111,
    240'b110000011111111110110110010100010101010101010101010101010101010101010101010100100101100010100001111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110111001111111111110101111,
    240'b110000011111111110110110010100010101010001010001010100000101001001010101010101010101010001010001011101111100011011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010010011111000011111111110101111,
    240'b110000011111111110110110010100000101011110000000100100010110100101010010010101010101010101010101010100010101011110000010110000011110111011111111111111111111111111111111111111111111111111111111111111001010100001011110111001001111111110101111,
    240'b110000011111111110110101010100001010100111111000111101011110001001101111010100100101010101010101010101010101010001010001010101010110110110010010101110011101001011100000111001111110011111010000100011100101010001011101111001011111111110101111,
    240'b110000011111111110110011011010011110111010100010011100011110000010110110010100100101010101010101010101010101010101010101010101000101001001010000010100010101011101100010011001110110011101011000010100010101001001011110111001011111111110110000,
    240'b110000011111111110110100010111111000100001011000010010001011110011001011010101000101010001010101010101010101010101010101010101010101010101010101010101010101010001010011010100100101001101010100010101010101001101011110111001011111111110110000,
    240'b110000011111111110110100010111011000010110001010100110111111000010100101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001011111111110110000,
    240'b110000011111111110110001011110101111100011110100111100001100000001100000010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001011111111110110000,
    240'b110000011111111110110001011111001110111010000100011010100101010101010010010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001011111111110110000,
    240'b101111101111111110110011011111001111011110111110101100101011011110000011010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110111001111111111110101011,
    240'b101101111111111111010001011101111101000111011100110111001101111010010100010011110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000100111101110101111101101111101110010101,
    240'b101100011111101111111100101010000110001101011110010111100101111001011100010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010110101111001100111111111110100010011111,
    240'b110001111101010011111111111111101110000011010110110101101101011011010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111110101011111111111111011100000011011000,
    240'b111011111100010011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110001001100110011110010,
    240'b111101111111010011000010101011111011110111000100110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111011100010110001110100111111011111110110,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule