module green_five(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100001111101111110100101010111001111010101010101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101011101010111010101110101011101010001001100110110000111011101111000111110001,
	240'b111100001111000111000100110100001110110011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110001110011111000111110000011110111011110001,
	240'b111011101100000011100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111100011111101110,
	240'b101111101101000011111111111101001010111010010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100011011000110010001100100011101011101011111100111111111100010010111001,
	240'b100011011111001111111110100110100100111101001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111101010011100000111000111110001110100011010111101110111000111111111101100110011011,
	240'b101000001111100011101101011001010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110110100111111001011101111111111001100000001111010111111101110100110101001,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010110011001100001101111101100011001110001111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010111011001111010111010111001111100011001110010111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110101110111111001111010011110011111001110001110011111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011000110001010000010110010101100001110101111110111111000110110011,
	240'b101100001111100111100110011000000101001101010011010100000100111101001111010100000101000001010001010100110101010101010101010101010101010101010101010101010101001001101110111100110111111001001110101110101010110101110001111110111111000110110011,
	240'b101100001111100111100110011000000100111101100100100101101010111110101100101000011000110001110010010111010101000101010001010101000101010101010101010101010101010001011001110011001110011011000111111101111000101001110001111110111111000110110011,
	240'b101100001111100111100110010111000111110011011111111111111111111111111111111111111111111011110110110110011010111001110111010101100101000101010101010101010101010101010011011010101011111111011000100110000101001001110101111110111111000110110011,
	240'b101100001111100111100011011110011110100011111111111111111111111111111111111111111111111111111111111111111111111111110101110001010111100101010010010100110101010101010101010100110101001101010101010100100101000001110101111110111111000110110011,
	240'b101100001111100011100010110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010101010010111010101000101010101010101010101010101010100010101010101000101110101111110111111000110110011,
	240'b101100001111011111101110111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000110110001010001010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111011011111001111101101111111111111111111111111111111111111111111111011110001011011011110111001101110011011100110111001101110011011100111000001101011101110011010100010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111011011111001111101111111111111111111111111111111111111111111111101000111100101011001010111000101110001011100010111000101110001011011011000011101110011100100011011110101000101010101010101010101000101110101111110111111000110110011,
	240'b101100001111011011110110111100111111111111111111111111111111111111111111111101000110111001001011010011100100111001001110010011100101000001010010010110011101010111111111110101100110000101010010010101010101000101110101111110111111000110110011,
	240'b101100001111011111110000111011001111111111111111111111111111111111111111111110011011010010100011101001011010010110100101101001111001000101010110010110011101010111111111111111111011100101010100010101000101000101110101111110111111000110110011,
	240'b101100001111100011100111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101011001010110001101010111111111111111111111101110001011010100000101000101110101111110111111000110110011,
	240'b101100001111100011100011110010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001101010001011001010110001101010111111111111111111111111111011110011000000100111101110101111110111111000110110011,
	240'b101100001111100011100000101001011111111111111111111111111111111111111111111111111111111111111101110011011001100110000110100001000111100001010101010110011101010111111111111111111111111111111111100111010100110001110101111110111111000110110011,
	240'b101100001111100111100010100000011111011011111111111111111111111111111111111111111111101010100001010110000100111001001110010011100100111101010001010101111101010011111111111111111111111111111111110111110101101101110011111110111111000110110011,
	240'b101100001111100111100100011001011101011111111111111111111111111111111111111111111011001101010010010100000101101101101100011011100110111001101101011100101101101111111111111111111111111111111111111111011000011101110000111110111111000110110011,
	240'b101100001111100111100110010110111010001111111111111111111111111111111111111100000110110001001110011100011101000111101101111011101110111011101110111011111111101111111111111111111111111111111111111111111011101101110011111110101111000110110011,
	240'b101100001111100111100110010111000110101111110000111111111111111111111111110100000101010101010101110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010010000011111110001111000110110011,
	240'b101100001111100111100110010111110101000010110101111111111111111111111111110000000101000101100100111010011111111111111111111111111111000011000001110000101111000011111111111111111111111111111111111111111111011110011110111101101111000110110011,
	240'b101100001111100111100110011000000101000001101101111011101111111111111111110010000101001101011011110110111111111111111111111111111100001001010001010111011101111111111111111111111111111111111111111111111111111110111101111101011111000110110011,
	240'b101100001111100111100110011000000101001101010001100111111111111111111111111001010110000101001111100011111111001111111111111010100111101101001100011100011111010111111111111111111111111111111111111111111111111111010110111101111111000110110011,
	240'b101100001111100111100110011000000101001101010011010110101100111011111111111111011001010101001110010100110111100010010100011011110101001001010000101011111111111111111111111111111111111111111111111111111111111111101011111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010100010110110111100100111111111110100101111000010011100100111001001110010011100100111110001011111101011111111111111111111111111111111111111111111111111111111111110111111111001111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101000001111101111011001111111111101010100110100110111001100100011100101010100011110011111111111111111111111111111111111111111111111111111111111111111111111100111111011111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010000100000011110100011111111111111111110111111100110111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111011111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010100000111010011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101111110011111000110110011,
	240'b101100001111100111100110011000000101001101010101010101000101010101010101010101010101000101100010101100001111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110000111101101111000110110011,
	240'b101100001111100111100110011000000101000101010011010110010101001101010011010101010101010101010011010100110111101011000011111101101111111111111111111111111111111111111111111111111111111111111111111111111100010001111010111110011111000110110011,
	240'b101100001111100111100110010111100101111010110110111000111011011101100001010100110101010101010101010101010101000101010110011110011011000011011010111101011111110111111111111111111111111111111010110001010110001001110010111110111111000110110011,
	240'b101100001111100111100101010111011011001011110000101101111110110110110100010100100101010101010101010101010101010101010100010100010101000101011101011100001000100110011100101001011010001010000000010110000100111001110101111110111111000110110011,
	240'b101100001111100111100101011001001100000110010101010001111001110111100010010111010101001101010101010101010101010101010101010101010101010101010011010100100101000001001111010011110100111101010001010101000101000101110101111110111111000110110011,
	240'b101100001111100111100110011000000101100001010111010101111011001111011011010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111100111100100011001101100000111100000111001011111010110010110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111100111100100011010011110001111001101101011001000010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111100111100100011010001110000110100010011010100111000001101000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110100111110111111000110110010,
	240'b100111011111100011101100011011111101110011111001111101001111011010111101010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111101111111111111101110100010100111,
	240'b100011011111000111111110101001000111010001111100011111010111110101101101010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011100101011110111111111111111101011110011010,
	240'b110000011100111011111111111110001011011010011001100110011001100110011011100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011101100111101100100011111110111111101100001010111100,
	240'b111011111100001011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101100100011101111,
	240'b111110011111001010111111110010011110010011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101001101111111000110110011001111100011111001,
	240'b111111111111100011100011101000101010000010110010101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100001001111010110111111111001111111111111110,
	240'b111100001111101111110100101010111001111010101010101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101011101010111010101110101011101010001001100110110000111011101111000111110001,
	240'b111100001111000111000100110100001110110011111000111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110001110011011000111110000011110111011110001,
	240'b111011101100000011100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111100011111101110,
	240'b101111101101000011111111111110011101011111001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110001101100010111000101110001101101110111111110111111111100010010111001,
	240'b100011011111001011111110110011001010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101001110000011100011111000111110001101011110111011011111111111101100110011011,
	240'b101000001111011111110110101100101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111010011111100011110111111111011101111110111101111111111110100110101001,
	240'b101100001111011111110011101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101100101011001010110000110111111110001010111000111111011111000110110011,
	240'b101100001111011111110011101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101100111011011100111100111110001010111000111111011111000110110011,
	240'b101100001111011111110011101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110111011111100111101001111001111100111010111001111111011111000110110011,
	240'b101100001111011111110011101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110101111110001100011010101000101011001010110010111010111111101111000110110011,
	240'b101100001111011111110011101011111010100110101001101010001010011110100111101001111010100010101000101010011010101010101010101010101010101010101010101010101010100010110111111110011011111010100111110111001101011010111000111111011111000110110011,
	240'b101100001111011111110011101011111010011110110010110010101101011111010101110100001100010110111001101011101010100010101000101010101010101010101010101010101010101010101100111001011111001011100011111110111100010010111000111111101111000110110011,
	240'b101100001111011111110011101011011011111011101111111111111111111111111111111111111111111011111010111011001101011010111011101010101010100010101010101010101010101010101001101101001101111111101100110010111010100010111010111111101111000110110011,
	240'b101100001111011111110001101111001111010011111111111111111111111111111111111111111111111111111111111111111111111111111010111000101011110010101001101010011010101010101010101010011010100110101010101010001010100010111010111111101111000110110011,
	240'b101100001111011111110001111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111010101101011101010100010101010101010101010101010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011011110111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001011010110101000101010101010101010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011011111101111110111111111111111111111111111111111111111111111111101111000011101101111011011110110111101101111011011110110111101101111100001110101110111001101010001010101010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011011111101111110111111111111111111111111111111111111111111111110101011110010101100101011011010110110101101101011011010111010101101101100001110110111110001101101111010100010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011011111011111110011111111111111111111111111111111111111111111110101011011010100101101001111010011110100111101001111010011110101000101010111110101011111111111010111011000010101001101010101010100010111010111111101111000110110011,
	240'b101100001111011011111000111101011111111111111111111111111111111111111111111111001101101011010001110100011101000111010001110100101100100010101010101011001110101011111111111111111101110010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011111110011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010101100101011001110101011111111111111111111110111000101101010001010100010111010111111101111000110110011,
	240'b101100001111011111110001111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110100110101100101011001110101011111111111111111111111111101110101011111010011110111010111111101111000110110011,
	240'b101100001111011111110000110100101111111111111111111111111111111111111111111111111111111111111110111001101100110011000010110000011011101110101010101011001110101011111111111111111111111111111111110011101010011010111010111111101111000110110011,
	240'b101100001111011111110001110000001111101011111111111111111111111111111111111111111111110011010000101010111010011110100110101001101010011110100111101010101110101011111111111111111111111111111111111011111010110110111001111111101111000110110011,
	240'b101100001111011111110010101100011110101111111111111111111111111111111111111111111101100110101000101010001010110110110110101101111011011110110110101110001110110111111111111111111111111111111111111111101100001110111000111111101111000110110011,
	240'b101100001111011111110011101011011101000111111111111111111111111111111111111110001011011010100110101110001110100011110110111101101111011011110111111101111111110111111111111111111111111111111111111111111101110110111001111111011111000110110011,
	240'b101100001111011111110011101011101011010111111000111111111111111111111111111001111010101010101010111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111000001111111001111000110110011,
	240'b101100001111011111110011101011111010100011011010111111111111111111111111110111111010100010110001111101001111111111111111111111111111100011100000111000001111100011111111111111111111111111111111111111111111101111001111111110111111000110110011,
	240'b101100001111011111110011101011111010100010110110111101101111111111111111111000111010100110101101111011011111111111111111111111111110000110101000101011101110111111111111111111111111111111111111111111111111111111011110111110111111000110110011,
	240'b101100001111011111110011101011111010100110101000110011111111111111111111111100101011000010100111110001111111100111111111111101001011110110100110101110001111101011111111111111111111111111111111111111111111111111101011111111001111000110110011,
	240'b101100001111011111110011101011111010100110101001101011011110011011111111111111101100101010100111101010011011110011001010101101111010100010101000110101111111111111111111111111111111111111111111111111111111111111110101111111011111000010110011,
	240'b101100001111011111110011101011111010100110101010101010001011011011110010111111111111010010111011101001111010011110100110101001111010011111000101111110101111111111111111111111111111111111111111111111111111111111111011111111101111000010110011,
	240'b101100001111011111110011101011111010100110101010101010101010100010111110111101101111111111110101110011011011011010110010101110011101001111111001111111111111111111111111111111111111111111111111111111111111111111111101111111111111000010110011,
	240'b101100001111011111110011101011111010100110101010101010101010101010101000101111111111001111111111111111111111011111110010111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111000010110011,
	240'b101100001111011111110011101011111010100110101010101010101010101010101010101010001011101011101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111111011111000110110011,
	240'b101100001111011111110011101011111010100110101010101010011010101010101010101010101010100010110001110101111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010111111110111111000110110011,
	240'b101100001111011111110011101011111010100010101001101011001010100110101001101010101010101010101001101010011011110111100001111110111111111111111111111111111111111111111111111111111111111111111111111111111110001010111101111111011111000110110011,
	240'b101100001111011111110011101011101010111011011010111100011101101110110000101010011010101010101010101010101010100010101010101111001101011111101100111110101111111011111111111111111111111111111100111000101011000010111001111111101111000110110011,
	240'b101100001111011111110011101011101101100011111000110110111111011011011001101010011010101010101010101010101010101010101010101010001010100010101110101110001100010011001101110100101101000010111111101011001010011110111010111111101111000110110011,
	240'b101100001111011111110010101100011110000011001010101000111100111011110000101011101010100110101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100010111010111111101111000110110011,
	240'b101100001111011111110011101011111010110010101011101010111101100111101101101011001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011111110010101100101110000011101111111100101111101011001011101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011111110010101101001111000111100110110101011100001010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111101111000110110011,
	240'b101100001111011111110010101101001111000011010001101101011011011110110100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111010111111101111000110110010,
	240'b100111011111011111110110101101111110111011111100111110011111101111011110101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011110111111111111111110100010100111,
	240'b100011011111000111111111110100011011100110111101101111101011111010110110101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010101111011111111111111101011110011010,
	240'b110000011100111011111111111110111101101011001100110011001100110011001101110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011111110001111111111111111101100001010111100,
	240'b111011111100001011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101100100011101111,
	240'b111110011111001010111111110010011110010011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101001101111111000110110011001111100011111001,
	240'b111111111111100011100011101000101010000010110010101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100001001111010110111111111001111111111111110,
	240'b111100001111101111110100101010111001111010101010101010111010101010101010101010101010101010101011101010111010101110101011101010111010101010101010101010101010101010101011101010111010101110101011101010001001100110110000111011101111000111110001,
	240'b111100001111000111000100110100001110110011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110001110011111000111110000011110111011110001,
	240'b111011101100000011100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111100011111101110,
	240'b101111101101000011111111111101001010111010010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100011011000110010001100100011101011101011111100111111111100010010111001,
	240'b100011011111001111111110100110100100111101001111010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111101010011100000111000111110001110100011010111101110111000111111111101100110011011,
	240'b101000001111100011101101011001010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110110100111111001011101111111111001100000001111010111111101110100110101001,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010110011001100001101111101100011001110001111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010111011001111010111010111001111100011001110010111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010110101110111111001111010011110011111001110001110011111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011000110001010000010110010101100001110101111110111111000110110011,
	240'b101100001111100111100110011000000101001101010011010100000100111101001111010100000101000001010001010100110101010101010101010101010101010101010101010101010101001001101110111100110111111001001110101110101010110101110001111110111111000110110011,
	240'b101100001111100111100110011000000100111101100100100101101010111110101100101000011000110001110010010111010101000101010001010101000101010101010101010101010101010001011001110011001110011011000111111101111000101001110001111110111111000110110011,
	240'b101100001111100111100110010111000111110011011111111111111111111111111111111111111111111011110110110110011010111001110111010101100101000101010101010101010101010101010011011010101011111111011000100110000101001001110101111110111111000110110011,
	240'b101100001111100111100011011110011110100011111111111111111111111111111111111111111111111111111111111111111111111111110101110001010111100101010010010100110101010101010101010100110101001101010101010100100101000001110101111110111111000110110011,
	240'b101100001111100011100010110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010101010010111010101000101010101010101010101010101010100010101010101000101110101111110111111000110110011,
	240'b101100001111011111101110111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000110110001010001010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111011011111001111101101111111111111111111111111111111111111111111111011110001011011011110111001101110011011100110111001101110011011100111000001101011101110011010100010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111011011111001111101111111111111111111111111111111111111111111111101000111100101011001010111000101110001011100010111000101110001011011011000011101110011100100011011110101000101010101010101010101000101110101111110111111000110110011,
	240'b101100001111011011110110111100111111111111111111111111111111111111111111111101000110111001001011010011100100111001001110010011100101000001010010010110011101010111111111110101100110000101010010010101010101000101110101111110111111000110110011,
	240'b101100001111011111110000111011001111111111111111111111111111111111111111111110011011010010100011101001011010010110100101101001111001000101010110010110011101010111111111111111111011100101010100010101000101000101110101111110111111000110110011,
	240'b101100001111100011100111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101011001010110001101010111111111111111111111101110001011010100000101000101110101111110111111000110110011,
	240'b101100001111100011100011110010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001101010001011001010110001101010111111111111111111111111111011110011000000100111101110101111110111111000110110011,
	240'b101100001111100011100000101001011111111111111111111111111111111111111111111111111111111111111101110011011001100110000110100001000111100001010101010110011101010111111111111111111111111111111111100111010100110001110101111110111111000110110011,
	240'b101100001111100111100010100000011111011011111111111111111111111111111111111111111111101010100001010110000100111001001110010011100100111101010001010101111101010011111111111111111111111111111111110111110101101101110011111110111111000110110011,
	240'b101100001111100111100100011001011101011111111111111111111111111111111111111111111011001101010010010100000101101101101100011011100110111001101101011100101101101111111111111111111111111111111111111111011000011101110000111110111111000110110011,
	240'b101100001111100111100110010110111010001111111111111111111111111111111111111100000110110001001110011100011101000111101101111011101110111011101110111011111111101111111111111111111111111111111111111111111011101101110011111110101111000110110011,
	240'b101100001111100111100110010111000110101111110000111111111111111111111111110100000101010101010101110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010010000011111110001111000110110011,
	240'b101100001111100111100110010111110101000010110101111111111111111111111111110000000101000101100100111010011111111111111111111111111111000011000001110000101111000011111111111111111111111111111111111111111111011110011110111101101111000110110011,
	240'b101100001111100111100110011000000101000001101101111011101111111111111111110010000101001101011011110110111111111111111111111111111100001001010001010111011101111111111111111111111111111111111111111111111111111110111101111101011111000110110011,
	240'b101100001111100111100110011000000101001101010001100111111111111111111111111001010110000101001111100011111111001111111111111010100111101101001100011100011111010111111111111111111111111111111111111111111111111111010110111101111111000110110011,
	240'b101100001111100111100110011000000101001101010011010110101100111011111111111111011001010101001110010100110111100010010100011011110101001001010000101011111111111111111111111111111111111111111111111111111111111111101011111110101111000110110011,
	240'b101100001111100111100110011000000101001101010101010100010110110111100100111111111110100101111000010011100100111001001110010011100100111110001011111101011111111111111111111111111111111111111111111111111111111111110111111111001111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101000001111101111011001111111111101010100110100110111001100100011100101010100011110011111111111111111111111111111111111111111111111111111111111111111111111100111111011111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010000100000011110100011111111111111111110111111100110111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111011111000110110011,
	240'b101100001111100111100110011000000101001101010101010101010101010101010101010100000111010011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101111110011111000110110011,
	240'b101100001111100111100110011000000101001101010101010101000101010101010101010101010101000101100010101100001111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110000111101101111000110110011,
	240'b101100001111100111100110011000000101000101010011010110010101001101010011010101010101010101010011010100110111101011000011111101101111111111111111111111111111111111111111111111111111111111111111111111111100010001111010111110011111000110110011,
	240'b101100001111100111100110010111100101111010110110111000111011011101100001010100110101010101010101010101010101000101010110011110011011000011011010111101011111110111111111111111111111111111111010110001010110001001110010111110111111000110110011,
	240'b101100001111100111100101010111011011001011110000101101111110110110110100010100100101010101010101010101010101010101010100010100010101000101011101011100001000100110011100101001011010001010000000010110000100111001110101111110111111000110110011,
	240'b101100001111100111100101011001001100000110010101010001111001110111100010010111010101001101010101010101010101010101010101010101010101010101010011010100100101000001001111010011110100111101010001010101000101000101110101111110111111000110110011,
	240'b101100001111100111100110011000000101100001010111010101111011001111011011010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111100111100100011001101100000111100000111001011111010110010110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111100111100100011010011110001111001101101011001000010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110101111110111111000110110011,
	240'b101100001111100111100100011010001110000110100010011010100111000001101000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110100111110111111000110110010,
	240'b100111011111100011101100011011111101110011111001111101001111011010111101010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111101111111111111101110100010100111,
	240'b100011011111000111111110101001000111010001111100011111010111110101101101010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011100101011110111111111111111101011110011010,
	240'b110000011100111011111111111110001011011010011001100110011001100110011011100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011101100111101100100011111110111111101100001010111100,
	240'b111011111100001011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101100100011101111,
	240'b111110011111001010111111110010011110010011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101001101111111000110110011001111100011111001,
	240'b111111111111100011100011101000101010000010110010101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100001001111010110111111111001111111111111110,
};
assign data = picture[addr];
endmodule