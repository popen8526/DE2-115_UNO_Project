module red_draw_two(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100001111001011101111110010011011010010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011010011000110111010011111001011110000,
	240'b111100011110001010111101110101101111000111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111000111010110101101111110000111110001,
	240'b111010101011100111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011100111101001,
	240'b101101001101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110111010,
	240'b100110001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110100101,
	240'b101010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111110111100101110111111101111111011111110111111110011011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111100110011000100110101001101001111010011110101001100111011001010111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111100010111110101111111111111111111111111111111111111111111011000110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111101100011100000111111111111111111111111111111111111111111101111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111110100011010001111111111111111111111111111111111111111111111011110000011110011111101100111100111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111100111000101111111101111111111111111111111111111111111111111110000001011101011001011110001001101010011111110111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111011001010111100011111111111111111111111111111111111111111110111101101101111111111111111011100110111101001111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111010110111000011111111111111111111111111111111111111111111011111100101111111111111111111110001111010101111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111101011110011101111111111111111111111111111111111111111111111001100010111111011111111111111011011000110111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111000110001111111110011111111111111111111111111111111111111111100110111101100111111111111111011000111111101101111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111110010011111001011111111111111111111111111111111111111111101111011011010111111111111111111010001111001111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111110110011101111011111111111111111111111111111111111111111111000111001010111111111111111111100101110100111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111011011100100011111010111111111111111111111111111111111111011111000001111110111111111111110100110010001111111011111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111101111011000011110000111100000110110010110001001011110111010011111111111111111111111111110001101111011011111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111101001111000110111100111011111111011011111111111111111111111111111111110101001110010011111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111011001111111111111111111111111111111111111111111001001101010011111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110100101111111111111111111111111111111111111111111101111100001011111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110100001100010111000110110001101100011011000110101111101101000111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111101101111011011110110111101101111011111111111011111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111,
	240'b101001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b100110011111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110100110,
	240'b101111101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010011000011,
	240'b111011101011101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001011100111101101,
	240'b111100111110100110111001110100011110110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110110111010010101101101110011111110011,
	240'b111100001111001111101111110010011011010110110110101101111011011010110110101101101011011010110110101101111011011110110111101101111011011110110110101101101011011010110110101101111011011110110111101101101011010111000110111010011111001111110000,
	240'b111100011110001010111100110101101111000111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111000111010110101101111110000111110001,
	240'b111010101011100111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011100111101001,
	240'b101101001101101011111111111100011010111010010000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100011111000110010001100100011111001000010010000100100001010110011101111111111111101101110111010,
	240'b100110001111101011111011100100000100111001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111010101110111110001110110010100100101000001010001010100000100111010001101111110101111101010100101,
	240'b101010001111111111100000010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110110001101111011011110110101011010101011001010100010101010101001101011011110111101111111110110011,
	240'b101011101111111111010100010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010010110111100011000110010100000111110000111101001010001010100100101001001011000110100101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110110100110100110100111001011001110000101000000101001101100100101000000001010011110100101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010010100111100010111110001001111010101010101100001110010110111101100001101101101110100101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010101111011110110110010000010100100101110011011011111111011111101011000110110100111111111110110111,
	240'b101011101111111111010101010110010101010001010100010100010101000001010000010100000101000101010011010101000101010101010101010101010101010101011100011000111010111011110100101100110110000101111111111000111100110001111010110100101111111110110111,
	240'b101011101111111111010101010110010101000101011010011111001001000010001110100001100111011001100101010101000101000001010010010101010101000010100111110011111001100011011000111111111000110101001011101000001000101101010010110100101111111110110111,
	240'b101011101111111111010101010101100111000011001011111110011111111111111111111111111111011011100100110001011001011101101001010100010100110110101000111011111110101011101000111010111000101001010001010101000101001101011000110100101111111110110111,
	240'b101011101111111111010010011011101101111111111111111111111111111111111111111111111111111111111111111111111111111111101001101011000110100101011011011010000110100101101001011010010101110001010100010101010101010001011000110100101111111110110111,
	240'b101011101111111111010010101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010010111010101010100111101010010010100100101010001010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111100010111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000100110010101010001010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111101110111110011111111111111111111111111111110111100101110111111101111111011111110111111110011011111100111111111111111111111111111111111101011001101101010100010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111110001111110101111111111111111111111111100110011000100110110001101100011011000110110011101000111001010111110101111111111111111111111111111111111011011011010110101000101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111101110111110001111111111111111111111111100010111110110110110101011000010101111101101001110001111011010110111011111111111111111111111111111111111111111110100110110000101010010010101010101010001011000110100101111111110110111,
	240'b101011101111111111101001111101111111111111111111111111111101100111011110100001110100101101010000010011010111001111011110110011011111111111111111111111111111111111111111111111111011101001010101010101000101010001011000110100101111111110110111,
	240'b101011101111111111100010111011101111111111111111111111111110100111010100100111010101000001010101010101000101001111000111110001101110011111101100111100111111111111111111111111111111110010010001010100000101010001011000110100101111111110110111,
	240'b101011101111111111011010110110111111111111111111111111111111100111001010110000010101001101010100010101010101000010100110110001011011111111010001110001101101010011111110111111111111111111100101011001100101000101011000110100101111111110110111,
	240'b101011101111111111010001101111101111111111111111111111111111111011001110110101010110001001010011010101010101000110000010110110011010110111001001111100001100111111101001111111111111111111111111101010110101000001011000110100101111111110110111,
	240'b101011101111111111001111100110101111111111111111111111111111111111011000110110110111110001010001010101010101001101100101110110100110011001001110100011111101111011010110111111111111111111111111111011000110100001010110110100101111111110110111,
	240'b101011101111111111010001011100111111000111111111111111111111111111101011110100011010000001010000010101010101010001010101110010101000101101001100010111001101010011001010111111111111111111111111111111111001111101010100110100101111111110110111,
	240'b101011101111111111010100010110111100110111111111111111111111111111111000110011001100000101010100010101010101010101010000101010001011010101001101010100101011101011001101111101101111111111111111111111111101011101011101110100011111111110110111,
	240'b101011101111111111010101010101001001000111111110111111111111111111111111110011001101100001100000010100010101010001001111100000001101001001010110010011111001100011010100111001111111111111111111111111111111011001111011110011101111111110110111,
	240'b101011101111111111010101010101110110000011100010111111111111111111111111110110101101110110011111010110010101101001010111011111111110110101101001010011100111010111011100110101001111111111111111111111111111111110100011110011011111111110110111,
	240'b101011101111111111010101010110010100111110011010111111111111111111111111111011011100100111110101110111011101100011011001111011001111111101111110010011010101110111010001110011001111111011111111111111111111111111000110110100001111111110110111,
	240'b101011101111111111010101010110010101001001011110110110001111111111111111111111111101111011000100110001111100010110110111101100111000100101010111010100110101001010111010110010111111011011111111111111111111111111100000110110101111111110110111,
	240'b101011101111111111010101010110010101010001010000100000001111011011111111111111111111111111111000111101001111000111000001110000110100111001010010010101010100111110010011110101101110010111111111111111111111111111110001111001001111111110110111,
	240'b101011101111111111010101010110010101010001010101010100101010011111111110111111111111111111111111111111111111111111010001111000011000001001010010010101010101000010001000111000101101010111111111111111111111111111111001111010111111111110110111,
	240'b101011101111111111010101010110010101010001010101010100110101100011000000111111111111111111111111111111111111111111100010110100111111000111001011110010001100100011100110111110001100001011111111111111111111111111111010111011101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101001101011111110001111111111111111111111111111111111111111101110100001100011111001010110010111100101111001001101111101101000111111111111111111111111111111011111100001111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010010011000001100000111111111111111111111111111111111111111101110111111101101111011011110110111101101111011111111111011111111111111111111111111111010111011011111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010100100101100110101011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111000001111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010001010001010100010100111101001111100000001101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001110011111111111110110111,
	240'b101011101111111111010101010110010101001101010100010101000110001001111011011110110111110001111100011001100101110010010110110101111111101111111111111111111111111111111111111111111111111111111111111111111101001101100110110100001111111110110111,
	240'b101011101111111111010101010110010101011001011000010100001000110111110111111100001111000011111010101100110100111001010000010111001000001010101111110101011110110011110101111110011111101011110000101110110110011001010101110100101111111110110111,
	240'b101011101111111111010100010100111001000110101110010011011000011011111111110110001000101110111001101000000101000101010101010101000101000001010001010110100110010101110111100000001000001001101110010101010101000101011000110100101111111110110111,
	240'b101011101111111111010101100001111101001011101001100100010101110110011011111100001100010001100011010101000101010101010101010101010101010101010101010101000101001101010001010100010101000101010010010101000101010001011000110100101111111110110111,
	240'b101011101111111111010101110000011111100011111100110110010101111101001101011111101110010011010001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111010100011000111011011111011001011001100101101001011100010100000110111011101011100111110101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111010100010101010111011010000110010011101000010011010010010111100100111011010001101101110101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111010101010110010101000101010001010100100111001011110011101101001001111011110100100100010101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101001011111111111100100010111110101001001010101010101010101001110011011111011011111001010111000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001011101111000101111111110110001,
	240'b100110011111011111111101100111010101001001010000010100000101000001001111011001110110110001010011010011110101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101001010011011111111001111011110100110,
	240'b101111101101001111111111111110001011111110100111101010001010100010101000101001011010010110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111011111011110111111111111101010011000011,
	240'b111011101011101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001011100111101101,
	240'b111100111110100110111001110100011110110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110110111010010101101101110011111110011,
	240'b111100001111001011101111110010011011010010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011010011000110111010011111001011110000,
	240'b111100011110001010111101110101101111000111110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111000111010110101101111110000111110001,
	240'b111010101011100111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011100111101001,
	240'b101101001101101011111111111100011010111010010000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100011111000110010001100100011111001000010010000100100001010110011101111111111111101101110111010,
	240'b100110001111101011111011100100000100111001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111010101110111110001110110010100100101000001010001010100000100111010001101111110101111101010100101,
	240'b101010001111111111100000010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011110110001101111011011110110101011010101011001010100010101010101001101011011110111101111111110110011,
	240'b101011101111111111010100010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010010110111100011000110010100000111110000111101001010001010100100101001001011000110100101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110110100110100110100111001011001110000101000000101001101100100101000000001010011110100101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000010010100111100010111110001001111010101010101100001110010110111101100001101101101110100101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010101111011110110110010000010100100101110011011011111111011111101011000110110100111111111110110111,
	240'b101011101111111111010101010110010101010001010100010100010101000001010000010100000101000101010011010101000101010101010101010101010101010101011100011000111010111011110100101100110110000101111111111000111100110001111010110100101111111110110111,
	240'b101011101111111111010101010110010101000101011010011111001001000010001110100001100111011001100101010101000101000001010010010101010101000010100111110011111001100011011000111111111000110101001011101000001000101101010010110100101111111110110111,
	240'b101011101111111111010101010101100111000011001011111110011111111111111111111111111111011011100100110001011001011101101001010100010100110110101000111011111110101011101000111010111000101001010001010101000101001101011000110100101111111110110111,
	240'b101011101111111111010010011011101101111111111111111111111111111111111111111111111111111111111111111111111111111111101001101011000110100101011011011010000110100101101001011010010101110001010100010101010101010001011000110100101111111110110111,
	240'b101011101111111111010010101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010010111010101010100111101010010010100100101010001010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111100010111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000100110010101010001010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111101110111110011111111111111111111111111111110111100101110111111101111111011111110111111110011011111100111111111111111111111111111111111101011001101101010100010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111110001111110101111111111111111111111111100110011000100110110001101100011011000110110011101000111001010111110101111111111111111111111111111111111011011011010110101000101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111101110111110001111111111111111111111111100010111110110110110101011000010101111101101001110001111011010110111011111111111111111111111111111111111111111110100110110000101010010010101010101010001011000110100101111111110110111,
	240'b101011101111111111101001111101111111111111111111111111111101100111011110100001110100101101010000010011010111001111011110110011011111111111111111111111111111111111111111111111111011101001010101010101000101010001011000110100101111111110110111,
	240'b101011101111111111100010111011101111111111111111111111111110100111010100100111010101000001010101010101000101001111000111110001101110011111101100111100111111111111111111111111111111110010010001010100000101010001011000110100101111111110110111,
	240'b101011101111111111011010110110111111111111111111111111111111100111001010110000010101001101010100010101010101000010100110110001011011111111010001110001101101010011111110111111111111111111100101011001100101000101011000110100101111111110110111,
	240'b101011101111111111010001101111101111111111111111111111111111111011001110110101010110001001010011010101010101000110000010110110011010110111001001111100001100111111101001111111111111111111111111101010110101000001011000110100101111111110110111,
	240'b101011101111111111001111100110101111111111111111111111111111111111011000110110110111110001010001010101010101001101100101110110100110011001001110100011111101111011010110111111111111111111111111111011000110100001010110110100101111111110110111,
	240'b101011101111111111010001011100111111000111111111111111111111111111101011110100011010000001010000010101010101010001010101110010101000101101001100010111001101010011001010111111111111111111111111111111111001111101010100110100101111111110110111,
	240'b101011101111111111010100010110111100110111111111111111111111111111111000110011001100000101010100010101010101010101010000101010001011010101001101010100101011101011001101111101101111111111111111111111111101011101011101110100011111111110110111,
	240'b101011101111111111010101010101001001000111111110111111111111111111111111110011001101100001100000010100010101010001001111100000001101001001010110010011111001100011010100111001111111111111111111111111111111011001111011110011101111111110110111,
	240'b101011101111111111010101010101110110000011100010111111111111111111111111110110101101110110011111010110010101101001010111011111111110110101101001010011100111010111011100110101001111111111111111111111111111111110100011110011011111111110110111,
	240'b101011101111111111010101010110010100111110011010111111111111111111111111111011011100100111110101110111011101100011011001111011001111111101111110010011010101110111010001110011001111111011111111111111111111111111000110110100001111111110110111,
	240'b101011101111111111010101010110010101001001011110110110001111111111111111111111111101111011000100110001111100010110110111101100111000100101010111010100110101001010111010110010111111011011111111111111111111111111100000110110101111111110110111,
	240'b101011101111111111010101010110010101010001010000100000001111011011111111111111111111111111111000111101001111000111000001110000110100111001010010010101010100111110010011110101101110010111111111111111111111111111110001111001001111111110110111,
	240'b101011101111111111010101010110010101010001010101010100101010011111111110111111111111111111111111111111111111111111010001111000011000001001010010010101010101000010001000111000101101010111111111111111111111111111111001111010111111111110110111,
	240'b101011101111111111010101010110010101010001010101010100110101100011000000111111111111111111111111111111111111111111100010110100111111000111001011110010001100100011100110111110001100001011111111111111111111111111111010111011101111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101001101011111110001111111111111111111111111111111111111111101110100001100011111001010110010111100101111001001101111101101000111111111111111111111111111111011111100001111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010010011000001100000111111111111111111111111111111111111111101110111111101101111011011110110111101101111011111111111011111111111111111111111111111010111011011111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010101010101010100100101100110101011111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111000001111111110110111,
	240'b101011101111111111010101010110010101010001010101010101010101010001010001010100010100111101001111100000001101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001110011111111111110110111,
	240'b101011101111111111010101010110010101001101010100010101000110001001111011011110110111110001111100011001100101110010010110110101111111101111111111111111111111111111111111111111111111111111111111111111111101001101100110110100001111111110110111,
	240'b101011101111111111010101010110010101011001011000010100001000110111110111111100001111000011111010101100110100111001010000010111001000001010101111110101011110110011110101111110011111101011110000101110110110011001010101110100101111111110110111,
	240'b101011101111111111010100010100111001000110101110010011011000011011111111110110001000101110111001101000000101000101010101010101000101000001010001010110100110010101110111100000001000001001101110010101010101000101011000110100101111111110110111,
	240'b101011101111111111010101100001111101001011101001100100010101110110011011111100001100010001100011010101000101010101010101010101010101010101010101010101000101001101010001010100010101000101010010010101000101010001011000110100101111111110110111,
	240'b101011101111111111010101110000011111100011111100110110010101111101001101011111101110010011010001011000010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111010100011000111011011111011001011001100101101001011100010100000110111011101011100111110101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111010100010101010111011010000110010011101000010011010010010111100100111011010001101101110101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101011101111111111010101010110010101000101010001010100100111001011110011101101001001111011110100100100010101000001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011000110100101111111110110111,
	240'b101001011111111111100100010111110101001001010101010101010101001110011011111011011111001010111000010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001011101111000101111111110110001,
	240'b100110011111011111111101100111010101001001010000010100000101000001001111011001110110110001010011010011110101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101001010011011111111001111011110100110,
	240'b101111101101001111111111111110001011111110100111101010001010100010101000101001011010010110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001111011111011110111111111111101010011000011,
	240'b111011101011101111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001011100111101101,
	240'b111100111110100110111001110100011110110111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110110111010010101101101110011111110011,
};
assign data = picture[addr];
endmodule