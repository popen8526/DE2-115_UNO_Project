module yellow_zero(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111110011111001111100110100111001000100110101001101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010111001001110001111111001001111111111101011,
	240'b111111001110001010111000110111001111010011111001111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111011011100110101111111110010011101111,
	240'b111101011011100011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111100000111011011,
	240'b101111101101011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110110010,
	240'b100111101111010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110,
	240'b101011001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000,
	240'b100111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101110,
	240'b101100011101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110101101,
	240'b111011011011100111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011111010000,
	240'b111111001101100010111011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110001101101010111101110,
	240'b111101011111111111100111101100111010101010101101101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101010101010101000110011111111011011100010,
	240'b111110011111001111100110100111001000100110101001101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010111001001110001111111001001111111111101011,
	240'b111111001110001010111000110111001111010011111010111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111011011100110101111111110010011101111,
	240'b111101011011100011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111100000111011011,
	240'b101111101101011011111111111101111101000111000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001011111110111101101111101100100111101111111111111110101110110010,
	240'b100111101111010011111110110010011010011010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101001101011010111001010101111101010011110111001111110001111111110101110,
	240'b101011001111111111110101101100011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101111001111010011111001111110101101000010101001111001011111111110110000,
	240'b101100101111111111110001101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111000001110101110110101110101001111010110110010110111111111111110110000,
	240'b101100101111111111110001101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101100111010101101001110100100101110101111010110111010110111111111111110110000,
	240'b101100101111111111110001101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101100111010101101001110100110101110101111010010111010110111111111111110110000,
	240'b101100101111111111110001101011111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101100111010101101001010100110101110011111010010111010110111111111111110110000,
	240'b101100101111111111110001101011111010100110101001101010001010100010101000101010001010100010101000101010011010101010101010101010101010101010101010101010101010101010101010111001111101111010100110110000111111011110110111110111111111111110110000,
	240'b101100101111111111110001101011111010011110110001110010011101011011010110110100101100100010111100101011111010100010101000101010011010101010101010101010101010101010101000110011001111101111100011111101011110010010101011111000001111111110110001,
	240'b101100101111111111110001101011011011110011101101111111111111111111111111111111111111111111111011111011111101101011000000101011001010100010101010101010101010101010101010101010111101000011101010110111101011010010101000111000011111111110110001,
	240'b101100101111111111101111101110111111001011111111111111111111111111111111111111111111111111111111111111111111111111111100111010001100001110101010101010001010101010101010101010101010100010101100101010011010100110101010111000011111111110110001,
	240'b101100101111111111101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011110101101001010100010101010101010101010101010101001101010101010101010101010111000011111111110110001,
	240'b101100101111111111110101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011100000010101000101010101010101010101010101010101010101010101010111000011111111110110001,
	240'b101100101111111111111001111111001111111111111111111111111111111111111111111111111111111111111111111111111111110111110100111100111111101111111111111111111111100011000111101010001010101010101010101010101010101010101010111000011111111110110001,
	240'b101100101111111111111001111111001111111111111111111111111111111111111111111111111111111111111111111010011100001010110011101100101011110011011111111111101111111111111010110001111010100010101010101010101010101010101010111000011111111110110000,
	240'b101100101111111111111000111111001111111111111111111111111111111111111111111111111111111111100010101011111010011110100111101001111010011110101010110100111111111011111111111110001011111010101000101010101010101010101010111000011111111110110000,
	240'b101100101111111111110110111110011111111111111111111111111111111111111111111111111111010010110101101001111010110111000001110001001011000010101000101011001110011011111111111111111110111110110010101010011010101010101010111000011111111110110000,
	240'b101100101111111111110011111100001111111111111111111111111111111111111111111111111101100110100111101010111101101011111110111111111110100110110001101001101100011011111111111111111111111111011101101010101010100110101010111000011111111110110000,
	240'b101100101111111111110000111001011111111111111111111111111111111111111111111111111100011010100101101111011111110111111111111111111111111111001101101001101011011111111010111111111111111111111100110000011010011110101010111000011111111110110000,
	240'b101100101111111111101110110101001111111111111111111111111111111111111111111111111100000010100101110001111111111111111111111111111111111111011001101001111011001111110110111111111111111111111111111010001010110010101001111000011111111110110001,
	240'b101100101111111111101111110000101111110011111111111111111111111111111111111111111100000010100101110001111111111111111111111111111111111111011001101001111011001111110101111111111111111111111111111111101100001010100111111000011111111110110001,
	240'b101100101111111111110000101100111110110111111111111111111111111111111111111111111100000010100101110001111111111111111111111111111111111111011001101001111011001111110101111111111111111111111111111111111110000110101001111000011111111110110001,
	240'b101100101111111111110001101011011101010011111111111111111111111111111111111111111100000010100101110001111111111111111111111111111111111111011001101001111011001111110101111111111111111111111111111111111111011110110101110111111111111110110001,
	240'b101100101111111111110001101011101011011111111001111111111111111111111111111111111100000010100101110001111111111111111111111111111111111111011001101001111011001111110101111111111111111111111111111111111111111111001001110111101111111110110001,
	240'b101100101111111111110001101011111010100011011110111111111111111111111111111111111100000010100101110001111111111111111111111111111111111111011001101001111011001111110101111111111111111111111111111111111111111111011110110111111111111110110000,
	240'b101100101111111111110001101011111010011110111001111110001111111111111111111111111100010010100101110000001111111011111111111111111111111111010010101001101011010111111000111111111111111111111111111111111111111111101101111001011111111110110000,
	240'b101100101111111111110001101011111010100110101000110101001111111111111111111111111101001110100111101011101110011111111111111111111111001110110111101001101100000111111110111111111111111111111111111111111111111111110111111010111111111110110000,
	240'b101100101111111111110001101011111010100110101001101011101110101011111111111111111110111110101111101001111011001011010010110101111011100110101000101010011101111111111111111111111111111111111111111111111111111111111100111100001111111110110000,
	240'b101100101111111111110001101011111010100110101010101010001011101011110101111111111111111111011000101010011010011110100111101001111010011110100111110010001111110011111111111111111111111111111111111111111111111111111101111101001111111110110000,
	240'b101100101111111111110001101011111010100110101010101010101010100011000100111110011111111111111110110110101011010110101010101010011011000111001111111110011111111111111111111111111111111111111111111111111111111111111101111101111111111110110000,
	240'b101100101111111111110001101011111010100110101010101010101010101010101000110001101111100111111111111111111111011011101000111001101111001011111111111111111111111111111111111111111111111111111111111111111111111111111101111101111111111110110001,
	240'b101100101111111111110001101011111010100110101010101010101010101010101010101010001100001011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100101111111110110001,
	240'b101100101111111111110001101011111010100110101010101010101010101010101010101010101010100010110111111000101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111001111111111110110001,
	240'b101100101111111111110001101011111010100110101000101010001010100010101010101010101010101010101000101010111100100011101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011110111111111111110110001,
	240'b101100101111111111110001101011111010100111000100110110101100100110101100101010011010101010101010101010011010100010110000110001111110010111110111111111111111111111111111111111111111111111111111111111001101010110101011111000001111111110110001,
	240'b101100101111111111110001101011011100100011111010111100001111101111010010101010011010101010101010101010101010101010101001101010001010101110110111110001111101011011100010111001101110100011011110110000101010101010101001111000011111111110110000,
	240'b101100101111111111110000101100001110101111011101101011001101001111110011101100001010100110101010101010101010101010101010101010101010101010101000101010001010100010101001101010111010110010101001101010001010101010101010111000011111111110110000,
	240'b101100101111111111110000101101001111000011001010101001001011111111110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101010101010101010111000011111111110110000,
	240'b101100101111111111110000101101001110111111001011101001011100000011110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111000011111111110110000,
	240'b101100101111111111110000101101001110111111001010101001001011111111110110101100111010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111000011111111110110000,
	240'b101100101111111111110000101100011110101111011100101010101101000111110011101100001010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111000011111111110110000,
	240'b101011111111111111110011101011101100101011111011111011111111101111010100101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111000111111111110110000,
	240'b100111111111011111111101101111111010011111000110110110111100101010101011101010001010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010011110110010111100111111111110101110,
	240'b101100011101111111111111111011111100000010110011101101001011001110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011101111100011111111111111000110101101,
	240'b111011011011100111110111111111111111110011110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111101011111111111111101100011111010000,
	240'b111111001101100010111011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110001101101010111101110,
	240'b111101011111111111100111101100111010101010101101101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101010101010101000110011111111011011100010,
	240'b111110011111001111100110100111001000100110101001101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010111001001110001111111001001111111111101011,
	240'b111111001110001010111000110111001111010111111011111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111110111111011011100110101111111110010011101111,
	240'b111101011011100011101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111100000111011011,
	240'b101111101101011011111111111001110111010001000011010000010100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100100001001000010010000100011111000111001001110110101111011001111111111111110101110110010,
	240'b100111101111010111111011010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000001111000000000000101101111010001111111110101110,
	240'b101011001111111111100000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101011101110111101100111100010111000100000000101100011111111110110000,
	240'b101100101111111111010011000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011100010000100110011111111110000000011000101000001111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000010111110000000000001100001110000100101111100111111111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000010111100100000000001100001101111100110000100111111111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000100111100000000000001011111101111100110001100111111111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101101111001101100000000010010111110011000100101101000001111111110110000,
	240'b101100101111111111010100000100000000000000010101010111011000010110000110011110010101100100110101000011110000000000000000000000000000000000000000000000000000000000000000011001101111001110101011111000001010111100000101101000111111111110110001,
	240'b101100101111111111010100000010110011011111001011111111111111111111111111111111111111111111110010110100001001001001000010000001110000000000000000000000000000000000000000000001100111001011000000100110110001110100000000101001001111111110110001,
	240'b101100101111111111001111001100111101011111111111111111111111111111111111111111111111111111111111111111111111111111110111101110100100101100000011000000000000000000000000000000000000000000000101000000000000000000000000101001001111111110110001,
	240'b101100101111111111010000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011110000111110000000000000000000000000000000000000000000000000000000000000000101001001111111110110001,
	240'b101100101111111111100010111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101000100001100000000000000000000000000000000000000000000000000000000101001001111111110110001,
	240'b101100101111111111101100111101111111111111111111111111111111111111111111111111111111111111111111111111111111101011011111110110111111010011111111111111111110101001010110000000000000000000000000000000000000000000000000101001001111111110110001,
	240'b101100101111111111101101111101111111111111111111111111111111111111111111111111111111111111111111101111000100101000011011000110010011011110011110111110111111111111110000010101100000000000000000000000000000000000000000101001001111111110110000,
	240'b101100101111111111101010111101101111111111111111111111111111111111111111111111111111111110101000000100000000000000000000000000000000000000000010011110111111110111111111111010100011110100000000000000000000000000000000101001001111111110110000,
	240'b101100101111111111100101111011011111111111111111111111111111111111111111111111111101111000011111000000000000100001000101010100000001001100000000000001111011011011111111111111111101000000011011000000000000000000000000101001001111111110110000,
	240'b101100101111111111011100110100111111111111111111111111111111111111111111111111111000110000000000000001011001000111111011111111111011101100010110000000000101010111111110111111111111111110011000000000100000000000000000101001001111111110110000,
	240'b101100101111111111010001101100011111111111111111111111111111111111111111111111110101010100000000001101111111011111111111111111111111111101101001000000000010011011101111111111111111111111110111010001100000000000000000101001001111111110110000,
	240'b101100101111111111001100011111111111111111111111111111111111111111111111111111110100001000000000010101101111111111111111111111111111111110001101000000000001110011100011111111111111111111111111101110100000100000000000101001001111111110110001,
	240'b101100101111111111001110010010011111010111111111111111111111111111111111111111110100000100000000010101101111111111111111111111111111111110001101000000000001110011100010111111111111111111111111111110110100100000000000101001001111111110110001,
	240'b101100101111111111010001000111001100100111111111111111111111111111111111111111110100000100000000010101101111111111111111111111111111111110001101000000000001110011100010111111111111111111111111111111111010011000000001101000111111111110110001,
	240'b101100101111111111010011000010100111111111111111111111111111111111111111111111110100000100000000010101101111111111111111111111111111111110001101000000000001110011100010111111111111111111111111111111111110011100100000101000001111111110110001,
	240'b101100101111111111010100000010110010100011101110111111111111111111111111111111110100000100000000010101101111111111111111111111111111111110001101000000000001110011100010111111111111111111111111111111111111111101011110100111011111111110110001,
	240'b101100101111111111010100000011110000000010011100111111111111111111111111111111110100000100000000010101101111111111111111111111111111111110001101000000000001110011100010111111111111111111111111111111111111111110011100100111111111111110110000,
	240'b101100101111111111010100000100000000000000101101111010111111111111111111111111110100111000000000010000111111110111111111111111111111111101110111000000000010001011101011111111111111111111111111111111111111111111001000101011111111111110110000,
	240'b101100101111111111010100000100000000000000000000011111101111111111111111111111110111110100000000000011011011011011111111111111111101101100100111000000000100011111111011111111111111111111111111111111111111111111100111110000101111111110110000,
	240'b101100101111111111010100000100000000000000000000000011101100000011111111111111111100111000010000000000000001100101111000100001110010111000000000000000001001111111111111111111111111111111111111111111111111111111110101110100111111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000011000011100010111111111111111110001001000000100000000000000000000000000000000000000000010110011111010111111111111111111111111111111111111111111111111111111000110111111111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000000000001001110111011101111111111111011100100010010010000000001000000000001100001110000111011101111111111111111111111111111111111111111111111111111111111111001111001101111111110110000,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000010101011110110111111111111111111110010010111001101101001101100011111111111111111111111111111111111111111111111111111111111111111111111111111010111001111111111110110001,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000100011111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110110001111111110110001,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000000000000101000101010001111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010101101011111111110110001,
	240'b101100101111111111010100000100000000000000000000000000000000000000000000000000000000000000000000000001010101100111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100011100111101111111110110001,
	240'b101100101111111111010100000011110000000001001110100100100101110100000110000000000000000000000000000000000000000000010010010110011011000011101000111111111111111111111111111111111111111111111111111101111000001000000101101000111111111110110001,
	240'b101100101111111111010100000010110101101011110001110100101111001001111001000000000000000000000000000000000000000000000000000000000000001100100111010110001000010110100111101101011011101010011110010010010000000100000000101001001111111110110000,
	240'b101100101111111111010010000100111100001010011010000011110111101111011010000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000010100000000000000000000000000000000101001001111111110110000,
	240'b101100101111111111010001000111101101000101100001000000000011111111100110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001001111111110110000,
	240'b101100101111111111010001000111101100111101100011000000000100000011100101000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001001111111110110000,
	240'b101100101111111111010001000111101101000001100001000000000011111111100110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001001111111110110000,
	240'b101100101111111111010010000101001100010010010101000010010111010111011100000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000111111111110110000,
	240'b101011111111111111011010000010110101111111110011110011101111010001111111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111110110000,
	240'b100111111111100011110111010000000000000001010100100101000110001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001110111001111111110101110,
	240'b101100011101111111111111110011100100010000011011000111100001110000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010011001110101011111111111111001010101101,
	240'b111011011011100111110111111111111111011011100010111000011110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000101110001011100010111000011110111111111111111111101100011111010000,
	240'b111111001101100010111011111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110001101101010111101110,
	240'b111101011111111111100111101100111010101010101101101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011101010101010101000110011111111011011100010,
};
assign data = picture[addr];
endmodule