module green_seven(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111100101111011011110010101101001010110010110101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101101010111110100111110111111111010011110010,
	240'b111011111111010011010111101111111101000111100110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111101011010111101110001001110110111110000,
	240'b111100011100111011001011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011100000111110001,
	240'b110010001100000111111101111111111101010110110010101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011011010110110101101101011011100100111111100111111111100100111001011,
	240'b100101101101111011111111110000110101101101001111010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001010011011011010111010001110011011100110111000110101110111111111110111110010010,
	240'b101000101110101111111101011111000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000110111001111010111110011111101101101100101110000111011011111101010011010,
	240'b101101111110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011001110110011100000001111010101100001110100101100110111000111111101010110000,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000101001111101000001001111011100101010011001100010111001001111101010110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111110101001110101010100000100111101011101111001011111101010110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101101101000110101010010100000101001101011101111001011111101010110001,
	240'b101110001110111011111000011011000101001001010100010100010100111101001111010100000101000101010011010101000101010101010101010101010101010101010101010101010101010101010101010100001001110011011011010110110101001001011101111001011111101010110001,
	240'b101110001110111011111000011011000100111101010110011110001001001110010010100010100111101001100101010101110101000001010010010101000101010101010101010101010101010101010101010100100110110011101010100000000100111101011101111001011111101010110001,
	240'b101110001110111011111000011010010110000010111101111101011111111111111111111111101111011011101011110010101001111101101110010101000101000101010101010101010101010101010101010101010101010010111110101001010101000001011101111001011111101010110001,
	240'b101110001110111011110111011100101100011011111111111111111111111111111111111111111111111111111111111111111111111111101111101111000111010001010010010100110101010101010101010101010101010001011100010111110101001101011101111001011111101010110001,
	240'b101110001110111011110011101010111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010101000010111000101000101010101010101010101010101010100010101000101001101011101111001011111101010110001,
	240'b101110001110111011111000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000110110101010001010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110110111111111111110011111111111111111111111111111111111111111111101101110110011101100111011001110110011101100111011001110110011101100111100001110000001111001010100000101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110110111111111111111001111111111111111111111111111111111111111101110110110010001100111011001110110011101100111011001110110011101100110011011001110001111101001011101110101000001010101010101010101001101011101111001011111101010110001,
	240'b101110001110110111111110111101011111111111111111111111111111111111111111101100010100111001010010010011100100110101001101010011010100111101010010010110001101100111111111111000010110101001010001010101010101001101011101111001011111101010110001,
	240'b101110001110110111111011111010101111111111111111111111111111111111111111101101110101000001011010100010011001001010010000100100101000000101010101010110101101101011111111111111111100101001011010010100110101001101011101111001011111101010110001,
	240'b101110001110111011110110110101111111111111111111111111111111111111111111110111000101110001010101110011101111111111111111111111111101001001010101010110001101101011111111111111111111111110011111010100000101001101011101111001011111101010110001,
	240'b101110001110111011110010101111111111111111111111111111111111111111111111111110111000000001001011100110011111111111111111111111111101001001010100010101111101101011111111111111111111111111101101011011010101000001011101111001011111101010110001,
	240'b101110001110111011110011100111101111110011111111111111111111111111111111111111111011010001001110011010101110111111111111111111111110111011000000110000011111000111111111111111111111111111111111101101100101000101011101111001011111101010110001,
	240'b101110001110111011110101100000001110101111111111111111111111111111111111111111111110010101100001010100011100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110110001011010111001011111101010110001,
	240'b101110001110111011111000011010111100010111111111111111111111111111111111111111111111110110001010010010111000111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111010010101011000111001011111101010110001,
	240'b101110001110111011111000011001111001000011111110111111111111111111111111111111111111111110111111010100000110010011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101100011111000111111101010110001,
	240'b101110001110111011111000011010100101111111100101111111111111111111111111111111111111111111101100011001110100111110111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000001111000011111101010110001,
	240'b101110001110111011111000011011000100110110100100111111111111111111111111111111111111111111111111100101000100101110000100111111001111111111111111111111111111111111111111111111111111111111111111111111111111111110100100110111111111101010110001,
	240'b101110001110111011111000011011000100111101100011111000111111111111111111111111111111111111111111110010100101001101011110111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111001000111000101111101010110001,
	240'b101110001110111011111000011011000101001001010000100100001111110011111111111111111111111111111111111100100110111101001101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111010001111100110110001,
	240'b101110001110111011111000011011000101001001010100010101101011111111111111111111111111111111111111111111111001111101001100011110111111100111111111111111111111111111111111111111111111111111111111111111111111111111101100111100101111100010110001,
	240'b101110001110111011111000011011000101001001010101010100100110010011011010111111111111111111111111111111111101001101010110010101111101011011111111111111111111111111111111111111111111111111111111111111111111111111110101111110001111011110110001,
	240'b101110001110111011111000011011000101001001010101010101010101000101110011111001001111111111111111111111111111011101111101010101011010101011111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111011110110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010000011101111110000111111111111111111111111111101000110110101110011011111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111011110110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010100010110110111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111100001111100010110001,
	240'b101110001110111011111000011011000101001001010100010101000101010101010101010101010101000101011110101010001111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111000101111101010110001,
	240'b101110001110111011111000011011000101001001011001010110000101010101010101010101010101010101010011010100100111011010111111111101001111111111111111111111111111111111111111111111111111111111111111111111111110011101110110111000101111101010110001,
	240'b101110001110111011111000011011000100111010001010101111110101101001010100010101010101010101010101010101010101000101010101011101101010110111011001111101101111111011111111111111111111111111111111110111110111110001011001111001011111101010110001,
	240'b101110001110111011111000011011000100111101110001111011010111101101010001010101010101010101010101010101010101010101010100010100010101000101011100011100101000101110100000101010111010110110010001011000100101000001011101111001011111101010110001,
	240'b101110001110111011111000011011000101000101010100110011001011000001010000010101010101010101010101010101010101010101010101010101010101010101010100010100100101000001010000010011110100111101010000010100110101001101011101111001011111101010110001,
	240'b101110001110111011111000011011000101001001010000100101011101111101011110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110111011111000011011000100110101001111011001111110100010000100010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110111011111000011010111000101001111001010011001100000010111011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110111011111000011010011101001110111100011001111010001011100110011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101001101110110011111011011101011100100011111011111100101111010111110100011011110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100100111011001111101010011110,
	240'b100100101110000111111111101101010111010101111111100000000111111101111011010101100100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101000010011101111111011111001110001100,
	240'b101111001100010111111111111111001011111010010111100101111001011110010111100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110101011011011110110111111111101000011000000,
	240'b111011101100011011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011110011101110,
	240'b111110011111011011000101110001101110000011110101111101111111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111001011111001,
	240'b111111111111110111101010101010101001110110110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100111010000110101001111100011111111111111111,
	240'b111100101111011011110010101101001010110010110101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101101010111110100111110111111111010011110010,
	240'b111011111111010011010111101111111101000111100110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111101011010111101110001001110110111110000,
	240'b111100011100111011001011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011100000111110001,
	240'b110010001100000111111101111111111110101011011000110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101101101011011010110110101101110010011111110111111111100100111001011,
	240'b100101101101111011111111111000011010110110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101001101101101011100110111001101110011011100011010110111111111110111110010010,
	240'b101000101110101011111110101111101010011110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101111111011101111101011111001111110101110110010111000111101111111100010011010,
	240'b101101111110111011111100101101011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100111011001110000010111101110110001111010010110011111100101111100010110000,
	240'b101110001110111011111100101101011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110100111110011110100111101110011101001010110001111100101111100010110001,
	240'b101110001110111011111100101101011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111010010111010101001111010011110101110111100101111100010110001,
	240'b101110001110111011111100101101011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111110100011010100101001111010100110101110111100101111100010110001,
	240'b101110001110111011111100101101011010100010101010101010001010011110100111101001111010100010101001101010101010101010101010101010101010101010101010101010101010101010101010101001111100110111101101101011011010100110101110111100101111100010110001,
	240'b101110001110111011111100101101011010011110101010101111001100100111001001110001011011110010110010101010111010011110101001101010101010101010101010101010101010101010101010101010011011010111110101101111111010011110101110111100101111100010110001,
	240'b101110001110111011111100101101001011000011011110111110101111111111111111111111101111101011110101111001011100111110110110101010011010100010101010101010101010101010101010101010101010101011011110110100101010011110101110111100101111100010110001,
	240'b101110001110111011111100101110001110001111111111111111111111111111111111111111111111111111111111111111111111111111110111110111011011101010101000101010011010101010101010101010101010101010101101101011111010100110101110111100101111100010110001,
	240'b101110001110111011111010110101011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011010100101011011010100010101010101010101010101010101001101010011010100110101110111100101111100010110001,
	240'b101110001110110111111101111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011011010101000101010101010101010101010101010101010100110101110111100101111100010110001,
	240'b101110001110110111111111111111001111111111111111111111111111111111111111111110111111010111110101111101011111010111110101111101011111010111110110111110001110111110111100101010001010101010101010101010101010100110101110111100101111100010110001,
	240'b101110001110110111111111111111011111111111111111111111111111111111111111110111011011000110110011101100111011001110110011101100111011001110110010101101101111000111110100101110111010100010101010101010101010100110101110111100101111100010110001,
	240'b101110001110110111111111111110101111111111111111111111111111111111111111110110001010011110101001101001111010011010100110101001101010011110101000101011001110110111111111111100001011010010101000101010101010100110101110111100101111100010110001,
	240'b101110001110110111111110111101011111111111111111111111111111111111111111110110111010100010101101110001001100100011000111110010001100000010101010101011001110110111111111111111111110010010101100101010011010100110101110111100101111100010110001,
	240'b101110001110110111111011111010111111111111111111111111111111111111111111111011011010110110101010111001111111111111111111111111111110100110101010101011001110110111111111111111111111111111001111101010001010100110101110111100101111100010110001,
	240'b101110001110111011111010110111111111111111111111111111111111111111111111111111011011111110100101110011001111111111111111111111111110100110101001101010111110110111111111111111111111111111110110101101101010100010101110111100101111100010110001,
	240'b101110001110111011111010110011101111110111111111111111111111111111111111111111111101101010100111101101011111011111111111111111111111011111100000111000001111100011111111111111111111111111111111110110111010100010101110111100101111100010110001,
	240'b101110001110111011111011101111111111010111111111111111111111111111111111111111111111001010110000101010001110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011011010101100111100101111100010110001,
	240'b101110001110111011111100101101011110001011111111111111111111111111111111111111111111111011000100101001011100011011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111101001010101100111100101111100010110001,
	240'b101110001110111011111100101100111100011111111111111111111111111111111111111111111111111111011111101010001011000111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010110001111100101111100010110001,
	240'b101110001110111011111100101101001010111111110010111111111111111111111111111111111111111111110101101100111010011111011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111000000111100001111100010110001,
	240'b101110001110111011111100101101011010011011010010111111111111111111111111111111111111111111111111110010101010010111000001111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111010010111100001111100010110001,
	240'b101110001110111011111100101101011010011110110001111100011111111111111111111111111111111111111111111001001010100110101110111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111100011111100010110001,
	240'b101110001110111011111100101101011010100010101000110010001111111011111111111111111111111111111111111110001011011110100110110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111101001111100010110001,
	240'b101110001110111011111100101101011010100010101010101010101101111111111111111111111111111111111111111111111100111110100101101111011111110011111111111111111111111111111111111111111111111111111111111111111111111111110110111110011111011110110001,
	240'b101110001110111011111100101101011010100010101010101010011011001011101100111111111111111111111111111111111110100110101011101010111110101111111111111111111111111111111111111111111111111111111111111111111111111111111010111111001111011110110001,
	240'b101110001110111011111100101101011010100010101010101010101010100010111001111100011111111111111111111111111111101110111110101010101101010011111111111111111111111111111111111111111111111111111111111111111111111111111100111111101111011110110001,
	240'b101110001110111011111100101101011010100010101010101010101010101010101000101110101111000011111111111111111111111111110100111011011111001111111111111111111111111111111111111111111111111111111111111111111111111111111100111111101111011110110001,
	240'b101110001110111011111100101101011010100010101010101010101010101010101010101010001011011011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111110001111011110110001,
	240'b101110001110111011111100101101011010100010101010101010101010101010101010101010101010100010101110110100111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111100011111100010110001,
	240'b101110001110111011111100101101011010100010101100101010111010101010101010101010101010101010101001101010001011101011011111111110011111111111111111111111111111111111111111111111111111111111111111111111111111001110111010111100011111100010110001,
	240'b101110001110111011111100101101011010011011000100110111111010110110101001101010101010101010101010101010101010100010101010101110101101011011101100111110101111111011111111111111111111111111111111111011111011111010101100111100101111100010110001,
	240'b101110001110111011111100101101011010011110111000111101101011110110101000101010101010101010101010101010101010101010101010101010001010100010101110101110001100010111010000110101011101011011001000101100011010011110101110111100101111100010110001,
	240'b101110001110111011111100101101011010100010101010111001101101100010101000101010101010101010101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100110101110111100101111100010110001,
	240'b101110001110111011111100101101011010100010100111110010101110111110101110101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101110111100101111100010110001,
	240'b101110001110111011111100101101011010011010100111101100111111001111000001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101110111100101111100010110001,
	240'b101110001110111011111100101101011100010010111100101001101101111111011101101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101110111100101111100010110001,
	240'b101110001110111011111100101101001110100111011110101100111101000011110011101100011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101110111100101111100010110001,
	240'b101001101110101111111110101110101110010011111101111110011111101011111001101101111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010110010111101101111100010011110,
	240'b100100101110000011111111110110101011101010111111101111111011111110111101101010111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011111001110111111111111001010001100,
	240'b101111001100010111111111111111101101111111001011110010111100101111001011110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011101101011111011111111111101000011000000,
	240'b111011101100011011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011110011101110,
	240'b111110011111011011000101110001101110000011110101111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111001011111001,
	240'b111111111111110111101010101010101001110110110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100111010000110101001111100011111111111111111,
	240'b111100101111011011110010101101001010110010110101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101101010111110100111110111111111010011110010,
	240'b111011111111010011010111101111111101000111100110111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111101011010111101110001001110110111110000,
	240'b111100011100111011001011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101011100000111110001,
	240'b110010001100000111111101111111111101010110110010101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011011010110110101101101011011100100111111100111111111100100111001011,
	240'b100101101101111011111111110000110101101101001111010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001010011011011010111010001110011011100110111000110101110111111111110111110010010,
	240'b101000101110101111111101011111000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100000110111001111010111110011111101101101100101110000111011011111101010011010,
	240'b101101111110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011001110110011100000001111010101100001110100101100110111000111111101010110000,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000101001111101000001001111011100101010011001100010111001001111101010110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100111110101001110101010100000100111101011101111001011111101010110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101101101000110101010010100000101001101011101111001011111101010110001,
	240'b101110001110111011111000011011000101001001010100010100010100111101001111010100000101000101010011010101000101010101010101010101010101010101010101010101010101010101010101010100001001110011011011010110110101001001011101111001011111101010110001,
	240'b101110001110111011111000011011000100111101010110011110001001001110010010100010100111101001100101010101110101000001010010010101000101010101010101010101010101010101010101010100100110110011101010100000000100111101011101111001011111101010110001,
	240'b101110001110111011111000011010010110000010111101111101011111111111111111111111101111011011101011110010101001111101101110010101000101000101010101010101010101010101010101010101010101010010111110101001010101000001011101111001011111101010110001,
	240'b101110001110111011110111011100101100011011111111111111111111111111111111111111111111111111111111111111111111111111101111101111000111010001010010010100110101010101010101010101010101010001011100010111110101001101011101111001011111101010110001,
	240'b101110001110111011110011101010111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000010101000010111000101000101010101010101010101010101010100010101000101001101011101111001011111101010110001,
	240'b101110001110111011111000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000110110101010001010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110110111111111111110011111111111111111111111111111111111111111111101101110110011101100111011001110110011101100111011001110110011101100111100001110000001111001010100000101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110110111111111111111001111111111111111111111111111111111111111101110110110010001100111011001110110011101100111011001110110011101100110011011001110001111101001011101110101000001010101010101010101001101011101111001011111101010110001,
	240'b101110001110110111111110111101011111111111111111111111111111111111111111101100010100111001010010010011100100110101001101010011010100111101010010010110001101100111111111111000010110101001010001010101010101001101011101111001011111101010110001,
	240'b101110001110110111111011111010101111111111111111111111111111111111111111101101110101000001011010100010011001001010010000100100101000000101010101010110101101101011111111111111111100101001011010010100110101001101011101111001011111101010110001,
	240'b101110001110111011110110110101111111111111111111111111111111111111111111110111000101110001010101110011101111111111111111111111111101001001010101010110001101101011111111111111111111111110011111010100000101001101011101111001011111101010110001,
	240'b101110001110111011110010101111111111111111111111111111111111111111111111111110111000000001001011100110011111111111111111111111111101001001010100010101111101101011111111111111111111111111101101011011010101000001011101111001011111101010110001,
	240'b101110001110111011110011100111101111110011111111111111111111111111111111111111111011010001001110011010101110111111111111111111111110111011000000110000011111000111111111111111111111111111111111101101100101000101011101111001011111101010110001,
	240'b101110001110111011110101100000001110101111111111111111111111111111111111111111111110010101100001010100011100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111100010110110001011010111001011111101010110001,
	240'b101110001110111011111000011010111100010111111111111111111111111111111111111111111111110110001010010010111000111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111010010101011000111001011111101010110001,
	240'b101110001110111011111000011001111001000011111110111111111111111111111111111111111111111110111111010100000110010011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101100011111000111111101010110001,
	240'b101110001110111011111000011010100101111111100101111111111111111111111111111111111111111111101100011001110100111110111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000001111000011111101010110001,
	240'b101110001110111011111000011011000100110110100100111111111111111111111111111111111111111111111111100101000100101110000100111111001111111111111111111111111111111111111111111111111111111111111111111111111111111110100100110111111111101010110001,
	240'b101110001110111011111000011011000100111101100011111000111111111111111111111111111111111111111111110010100101001101011110111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111001000111000101111101010110001,
	240'b101110001110111011111000011011000101001001010000100100001111110011111111111111111111111111111111111100100110111101001101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111010001111100110110001,
	240'b101110001110111011111000011011000101001001010100010101101011111111111111111111111111111111111111111111111001111101001100011110111111100111111111111111111111111111111111111111111111111111111111111111111111111111101100111100101111100010110001,
	240'b101110001110111011111000011011000101001001010101010100100110010011011010111111111111111111111111111111111101001101010110010101111101011011111111111111111111111111111111111111111111111111111111111111111111111111110101111110001111011110110001,
	240'b101110001110111011111000011011000101001001010101010101010101000101110011111001001111111111111111111111111111011101111101010101011010101011111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111011110110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010000011101111110000111111111111111111111111111101000110110101110011011111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111011110110001,
	240'b101110001110111011111000011011000101001001010101010101010101010101010101010100010110110111010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111100001111100010110001,
	240'b101110001110111011111000011011000101001001010100010101000101010101010101010101010101000101011110101010001111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111000101111101010110001,
	240'b101110001110111011111000011011000101001001011001010110000101010101010101010101010101010101010011010100100111011010111111111101001111111111111111111111111111111111111111111111111111111111111111111111111110011101110110111000101111101010110001,
	240'b101110001110111011111000011011000100111010001010101111110101101001010100010101010101010101010101010101010101000101010101011101101010110111011001111101101111111011111111111111111111111111111111110111110111110001011001111001011111101010110001,
	240'b101110001110111011111000011011000100111101110001111011010111101101010001010101010101010101010101010101010101010101010100010100010101000101011100011100101000101110100000101010111010110110010001011000100101000001011101111001011111101010110001,
	240'b101110001110111011111000011011000101000101010100110011001011000001010000010101010101010101010101010101010101010101010101010101010101010101010100010100100101000001010000010011110100111101010000010100110101001101011101111001011111101010110001,
	240'b101110001110111011111000011011000101001001010000100101011101111101011110010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110111011111000011011000100110101001111011001111110100010000100010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110111011111000011010111000101001111001010011001100000010111011010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101110001110111011111000011010011101001110111100011001111010001011100110011000100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101111001011111101010110001,
	240'b101001101110110011111011011101011100100011111011111100101111010111110100011011110101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100100111011001111101010011110,
	240'b100100101110000111111111101101010111010101111111100000000111111101111011010101100100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101000010011101111111011111001110001100,
	240'b101111001100010111111111111111001011111010010111100101111001011110010111100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110101011011011110110111111111101000011000000,
	240'b111011101100011011010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011110011101110,
	240'b111110011111011011000101110001101110000011110101111101111111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101110010111001100110000111111001011111001,
	240'b111111111111110111101010101010101001110110110001101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100111010000110101001111100011111111111111111,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule