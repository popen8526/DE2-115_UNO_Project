module blue_one(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111110111111001011011110100111101010011011000001110000111100001111000011110000111100001011000010110000101100001011000010110000111100001111000011110000111100001111000010110000101100001011000011101111101001111110110001111101111111111111111001,
	240'b111111001110101010111100110010001110001011100100111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001110000011000100110011111111110111111010,
	240'b111110111011110011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001101001011111100,
	240'b110011011101000111111111111101111100000010100100101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100000101000111100110011111101111111111100100011001101,
	240'b101001001111001111111101100111010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101101111011011110101010010111010111111111110010010011100,
	240'b101011101111111111101000011000010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011000010111100010111110101110101111110101111001110101101,
	240'b101101001111111111011010010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011000110111100001011111101101111111100011111010010110111,
	240'b101101001111111111011010010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011001000101110000111100001110010111100011111010010110111,
	240'b101101001111111111011010010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011001001101100110100110001101110111100101111010010110111,
	240'b101101001111111111011010010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011001001101101000100111001101110111100101111010010110111,
	240'b101101011111111111011010010111000101010001010011010100000101000001010000010100000101000101010011010101000101010101010101010101010101010101010101010101010101010101010101010101000101010011001001101101000100111001101110111100101111010010110111,
	240'b101101011111111111011010010111000101000001011101100000101001100010010110100010110111101001100110010101010101000001010010010101010101010101010101010101010101010101010101010101000101010011001011101101100100111001101110111100101111010010110111,
	240'b101101011111111111011010010110000111011111010100111111001111111111111111111111111111011111101000110010001001101101101100010100100101001001010101010101010101010101010101010101000101010010110111101001010100111001101110111100101111010010110111,
	240'b101101011111111111010111011101001110010011111111111111111111111111111111111111111111111111111111111111111111111111101100101100100110110001010001010101000101010101010101010101010101010101011110010111000101001001101110111100101111010010110111,
	240'b101101011111111111011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110011010010101110101001001010101010101010101010101010100010101000101001001101110111100101111010010110111,
	240'b101101011111111111100111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111110110001001010001010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111110000111110011111111111111111111111111111111111111111111111111111111111111111111111111111010011101010111011101111111111111111111111111101010001101010010100010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111110001111110011111111111111111111111111111111111111111111111111111111111111111111111111010101001100000011001111100000011111111111111111111111111011000011010010101000101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111101111111110011111111111111111111111111111111111111111111111111111111111111111111111111010000001001110010100000101111111001101111111111111111111111111110011110101111001010011010101010101001001101110111100101111010010110111,
	240'b101101001111111111101010111101011111111111111111111111111111111111111111111111111111111111111111111111111010000101010000010101010100111101101001111001001111111111111111111111111011001101010100010101000101001001101110111100101111010010110111,
	240'b101101001111111111100011111001111111111111111111111111111111111111111111111111111111111111111111111111111010000101001110011010110111010101010001110010111111111111111111111111111111101010001000010100000101001001101110111100101111010010110111,
	240'b101101011111111111011011110100101111111111111111111111111111111111111111111111111111111111111111111111111010000101001100011110111101110001110011110010001111111111111111111111111111111111011101011000000101000001101110111100101111010010110111,
	240'b101101011111111111010101101100011111111111111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111101111011100110111001111111111111111111111111111111111111111100111010100110101101110111100101111010010110111,
	240'b101101011111111111010110100011001111110011111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111000000101110001101100111100101111010010110111,
	240'b101101011111111111011000011010011110010011111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111101000101001101001111100101111010010110111,
	240'b101101011111111111011010010110011011010111111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111100000001101101111100101111010010110111,
	240'b101101011111111111011010010110000111100111111000111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111110100001111111111100001111010010110111,
	240'b101101001111111111011010010110110101010111000111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111101010011101111011011111010010110111,
	240'b101101001111111111011010010111000100111101111100111101111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111111110111110111011011111010010110111,
	240'b101101001111111111011010010111000101001101010011101101001111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111011010111011111111001110110111,
	240'b101101001111111111011010010111000101010001010010011001001101111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111101011111100101111001110110111,
	240'b101101001111111111011010010111000101010001010101010100010111110011110000111111111111111111111111111111111010000001001011011101101111011111111111111111111111111111111111111111111111111111111111111111111111111111110001111101011111001110110111,
	240'b101101011111111111011010010111000101010001010101010101010101000010001111111101101111111111111111111111111010010001010010011111001111011111111111111111111111111111111111111111111111111111111111111111111111111111110011111101111111001110110111,
	240'b101101011111111111011010010111000101010001010101010101010101010101010001100100111111010111111111111111111110100011010011110111101111110111111111111111111111111111111111111111111111111111111111111111111111111111110100111101111111001110110111,
	240'b101101011111111111011010010111000101010001010101010101010101010101010100010100011000010111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111100101111001110110111,
	240'b101101011111111111011010010111000101010001010100010101000101010101010101010101010101000001101111110001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111011101111010010110111,
	240'b101101011111111111011010010111000101010001011000010101110101010101010101010101010101010101010001010110011001000011011000111111011111111111111111111111111111111111111111111111111111111111111111111111111101101101111110111100001111010010110111,
	240'b101101011111111111011010010110110101010110101110100100000101000101010101010101010101010101010101010101000101000001011101100010101100001011101001111110111111111111111111111111111111111111111111110111000111001101101010111100101111010010110111,
	240'b101101001111111111011010010110110101011011010110101010100100111101010101010101010101010101010101010101010101010101010011010100000101010101100110100000101001101010101101101101111011010110010110011000110100111001101110111100101111010010110111,
	240'b101101001111111111011010010110110101011011010011101010000100111101010101010101010101010101010101010101010101010101010101010101010101010001010011010100000101000001010010010100110101001001010000010100110101001001101110111100101111010010110111,
	240'b101101001111111111011010010110110101011011010011101010000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111011010010110100101010011010011101010000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111011001011001000110111011010010101010000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101011111111111011000011011011100111111101100101001100100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101100001111111111100011010111101010110011111111101001010100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101111111010010110001,
	240'b101000111111011111111011100010100101001110001010011011110100111001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000010101000111111111110100110011100,
	240'b110000111101100111111111111011011010000110000010100001101000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011011000011110111111111111100110011000000,
	240'b111101111011100111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011100101111111000,
	240'b111110001110101110111111110111001110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011010001101111101110111111111000,
	240'b111100111111111111110001101000001000111110101010101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101001111000100010101000111010111111000011110101,
	240'b111110111111001011011110100111101010011011000001110000111100001111000011110000111100001011000010110000101100001011000010110000111100001111000011110000111100001111000010110000101100001011000011101111101001111110110001111101111111111111111001,
	240'b111111001110101010111100110010001110001011100100111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001001110000011000100110011111111110111111010,
	240'b111110111011110011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001101001011111100,
	240'b110011011101000111111111111101111100000010100100101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100000101000111100110011111101111111111100100011001101,
	240'b101001001111001111111101100111010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101101111011011110101010010111010111111111110010010011100,
	240'b101011101111111111101000011000010101001001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011000010111100010111110101110101111110101111001110101101,
	240'b101101001111111111011010010110110101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011000110111100001011111101101111111100011111010010110111,
	240'b101101001111111111011010010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011001000101110000111100001110010111100011111010010110111,
	240'b101101001111111111011010010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011001001101100110100110001101110111100101111010010110111,
	240'b101101001111111111011010010111000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010011001001101101000100111001101110111100101111010010110111,
	240'b101101011111111111011010010111000101010001010011010100000101000001010000010100000101000101010011010101000101010101010101010101010101010101010101010101010101010101010101010101000101010011001001101101000100111001101110111100101111010010110111,
	240'b101101011111111111011010010111000101000001011101100000101001100010010110100010110111101001100110010101010101000001010010010101010101010101010101010101010101010101010101010101000101010011001011101101100100111001101110111100101111010010110111,
	240'b101101011111111111011010010110000111011111010100111111001111111111111111111111111111011111101000110010001001101101101100010100100101001001010101010101010101010101010101010101000101010010110111101001010100111001101110111100101111010010110111,
	240'b101101011111111111010111011101001110010011111111111111111111111111111111111111111111111111111111111111111111111111101100101100100110110001010001010101000101010101010101010101010101010101011110010111000101001001101110111100101111010010110111,
	240'b101101011111111111011000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100110011010010101110101001001010101010101010101010101010100010101000101001001101110111100101111010010110111,
	240'b101101011111111111100111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111110110001001010001010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111110000111110011111111111111111111111111111111111111111111111111111111111111111111111111111010011101010111011101111111111111111111111111101010001101010010100010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111110001111110011111111111111111111111111111111111111111111111111111111111111111111111111010101001100000011001111100000011111111111111111111111111011000011010010101000101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111101111111110011111111111111111111111111111111111111111111111111111111111111111111111111010000001001110010100000101111111001101111111111111111111111111110011110101111001010011010101010101001001101110111100101111010010110111,
	240'b101101001111111111101010111101011111111111111111111111111111111111111111111111111111111111111111111111111010000101010000010101010100111101101001111001001111111111111111111111111011001101010100010101000101001001101110111100101111010010110111,
	240'b101101001111111111100011111001111111111111111111111111111111111111111111111111111111111111111111111111111010000101001110011010110111010101010001110010111111111111111111111111111111101010001000010100000101001001101110111100101111010010110111,
	240'b101101011111111111011011110100101111111111111111111111111111111111111111111111111111111111111111111111111010000101001100011110111101110001110011110010001111111111111111111111111111111111011101011000000101000001101110111100101111010010110111,
	240'b101101011111111111010101101100011111111111111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111101111011100110111001111111111111111111111111111111111111111100111010100110101101110111100101111010010110111,
	240'b101101011111111111010110100011001111110011111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111000000101110001101100111100101111010010110111,
	240'b101101011111111111011000011010011110010011111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111101000101001101001111100101111010010110111,
	240'b101101011111111111011010010110011011010111111111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111100000001101101111100101111010010110111,
	240'b101101011111111111011010010110000111100111111000111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111110100001111111111100001111010010110111,
	240'b101101001111111111011010010110110101010111000111111111111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111101010011101111011011111010010110111,
	240'b101101001111111111011010010111000100111101111100111101111111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111111110111110111011011111010010110111,
	240'b101101001111111111011010010111000101001101010011101101001111111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111011010111011111111001110110111,
	240'b101101001111111111011010010111000101010001010010011001001101111111111111111111111111111111111111111111111010000101001100011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111101011111100101111001110110111,
	240'b101101001111111111011010010111000101010001010101010100010111110011110000111111111111111111111111111111111010000001001011011101101111011111111111111111111111111111111111111111111111111111111111111111111111111111110001111101011111001110110111,
	240'b101101011111111111011010010111000101010001010101010101010101000010001111111101101111111111111111111111111010010001010010011111001111011111111111111111111111111111111111111111111111111111111111111111111111111111110011111101111111001110110111,
	240'b101101011111111111011010010111000101010001010101010101010101010101010001100100111111010111111111111111111110100011010011110111101111110111111111111111111111111111111111111111111111111111111111111111111111111111110100111101111111001110110111,
	240'b101101011111111111011010010111000101010001010101010101010101010101010100010100011000010111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010111100101111001110110111,
	240'b101101011111111111011010010111000101010001010100010101000101010101010101010101010101000001101111110001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111011101111010010110111,
	240'b101101011111111111011010010111000101010001011000010101110101010101010101010101010101010101010001010110011001000011011000111111011111111111111111111111111111111111111111111111111111111111111111111111111101101101111110111100001111010010110111,
	240'b101101011111111111011010010110110101010110101110100100000101000101010101010101010101010101010101010101000101000001011101100010101100001011101001111110111111111111111111111111111111111111111111110111000111001101101010111100101111010010110111,
	240'b101101001111111111011010010110110101011011010110101010100100111101010101010101010101010101010101010101010101010101010011010100000101010101100110100000101001101010101101101101111011010110010110011000110100111001101110111100101111010010110111,
	240'b101101001111111111011010010110110101011011010011101010000100111101010101010101010101010101010101010101010101010101010101010101010101010001010011010100000101000001010010010100110101001001010000010100110101001001101110111100101111010010110111,
	240'b101101001111111111011010010110110101011011010011101010000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111011010010110100101010011010011101010000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101001111111111011001011001000110111011010010101010000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101101011111111111011000011011011100111111101100101001100100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101110111100101111010010110111,
	240'b101100001111111111100011010111101010110011111111101001010100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110011111101111111010010110001,
	240'b101000111111011111111011100010100101001110001010011011110100111001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000010101000111111111110100110011100,
	240'b110000111101100111111111111011011010000110000010100001101000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011011000011110111111111111100110011000000,
	240'b111101111011100111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011100101111111000,
	240'b111110001110101110111111110111001110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011010001101111101110111111111000,
	240'b111100111111111111110001101000001000111110101010101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101001111000100010101000111010111111000011110101,
	240'b111110111111001011011110100111101010011011000001110000111100001111000011110000111100001011000010110000101100001011000010110000111100001111000011110000111100001111000010110000101100001011000011101111101001111110110001111101111111111111111001,
	240'b111111001110101010111100110010001110001011100100111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111001011110010111100101111000111101111111000100110011111111110111111010,
	240'b111110111011110011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100001101001011111100,
	240'b110011011101000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100011001101,
	240'b101001001111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010010011100,
	240'b101011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010101101,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110111,
	240'b101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010110001,
	240'b101000111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010011100,
	240'b110000111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011000000,
	240'b111101111011100111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011100101111111000,
	240'b111110001110101110111111110111001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111010001101111101110111111111000,
	240'b111100111111111111110001101000001000111110101010101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101101101001111000100010101000111010111111000011110101,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule