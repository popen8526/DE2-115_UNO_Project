module green_four(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111100101111110011100111101011001010111110110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011010110010101011111001101111010011110011,
	240'b111100001111100011001101110000011101011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111101001010111011110010011110111111110000,
	240'b111100011100011011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001100100011110011,
	240'b110010101100101111111111111110111100101010110001101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001010111010101110101100101101001111111111111111101100001011001010,
	240'b100101111111001111111110101010000101010001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010110101101100010010011100101101010111110111111111110001010011001,
	240'b100111101111111011101011011001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011010110011001011010101100100111101110110111110101111001110100100,
	240'b101011101111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000111000011101101011111010100111001101010111100011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011011001001001111001010101111100100111101101010111100011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100011011110100110001011111010010110101101100111111100011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100011001110100001100001110100111010100101100110111100011111110010101111,
	240'b101011111111111011011110010111010101010001010100010100010100111101001111010100000101000101010011010101000101010101010101010101010101010101010101010101010101001101100001110101111111101011010110111100011101100001101110111100001111110010101111,
	240'b101011111111111011011110010111010101000001011011100000001001010010010001100010000111011001100010010101010101000001010011010101010101010101010101010101010101001101011110110011001111101011000100101111101010000101101110111100001111110010101111,
	240'b101011111111111011011110010110010111000011001110111110011111111111111111111111011111010011100111110000111001011001100111010100100101001001010101010101010101010101010000100000101101011001011000010011100100111001101011111100011111110010101111,
	240'b101011111111111011011011011100011101111111111111111111111111111111111111111111111111111111111111111111111111111111101000101011110110101001010001010101000101010101010101010110010110000101010110010101010101001001101011111100011111110010101111,
	240'b101011111111111011011011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010011001010101110101001001010101010101000101001101010101010101010101001001101011111100011111110010101111,
	240'b101011111111110011100111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111100110001101010001010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111101111110100111101101111111111111111111111111111111111111111111111111111111111111111111111011110110111101011111101101111111111111111111111111101010101101010010100010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111101111110101111101111111111111111111111111111111111111111111111111111111111111111111111110111001000001011111100101001111110111111111111111111111111111011001011010010101000101010101010101010101001001101011111100011111110010101111,
	240'b101011111111101111110010111101001111111111111111111111111111111111111111111111111111111111111111111111111011111001001111010110111101101111111111111111111111111111111111110100000101111101010011010101010101001001101011111100011111110010101111,
	240'b101011111111110011101100111100001111111111111111111111111111111111111111111111111111111111111111111111111111001101110001010011001001110011111111111111111111111111111111111111111011011001010100010101000101001001101011111100011111110010101111,
	240'b101011111111110111100011111001101111111111111111111111111111111111111111111111111111111111111111111111111111111110101110010011100110010111101000111111111111111111111111111111111111101010001011010100000101001001101011111100011111110010101111,
	240'b101011111111110111011101110100001111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011001010100111010101110111111111111111111111111111111111111111111011111011000010101000001101011111100011111110010101111,
	240'b101011111111111011011001101011101111111111111111111111111111111111111111111111111111111111110100101000101001000111010011100111110100110001110010111100111111111111111111111111111111111111111111101000100100110101101011111100011111110010101111,
	240'b101011111111111011011001100010011111101111111111111111111111111111111111111111111111111111101110011001100100101010110110111000000101110001010010110000001111111111111111111111111111111111111111111000110101111101101000111100011111110010101111,
	240'b101011111111111011011100011001111110000111111111111111111111111111111111111111111111111111101110011010100100111110110101111111111000101101001011100000001111101011111111111111111111111111111111111111101000111101100110111100011111110010101111,
	240'b101011111111111011011110010110011011000011111111111111111111111111111111111111111111111111101110011010100100111110110100111111111100101101010101010101111101000111111111111111111111111111111111111111111100010101101010111100001111110010101111,
	240'b101011111111111011011110010110010111010111110110111111111111111111111111111111111111111111110010011010110100111110110111111111111111110001111110010011001001000111111101111111111111111111111111111111111110101101111111111011101111110010101111,
	240'b101011111111111011011110010111000101001111000010111111111111111111111111111111111110101111000000011001000101000110011000110100001101000110010100010100000110000011100100111111111111111111111111111111111111110010011110111011001111110010101111,
	240'b101011111111111011011110010111010100111101110111111101011111111111111111111111111011011101010011010101010101010101010111010110000101100001011000010101000101011011010100111111111111111111111111111111111111111111000000111011001111110010101111,
	240'b101011111111111011011110010111010101001101010010101011011111111111111111111111111011010001001100010101000101010101010011010100010101000101010001010100010101010011010100111111111111111111111111111111111111111111011001111100001111110010101111,
	240'b101011111111111011011110010111010101010001010011010111111101100011111111111111111101111010100100011000000101001010001000101100011011000010110000101011111011000011101011111111111111111111111111111111111111111111101101111101001111101110101111,
	240'b101011111111111011011110010111010101010001010101010100010111011011101100111111111111111111110010011010010100110110110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101111111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101000010000110111100011111111111101111011100100101100010111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110001111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010001100010101110111011111111111000011101101111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110001111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010100000111110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111101001111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101010001010101010101010101000101100111101110001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111000111011011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101100101010110010101010101010101010010010101001000000111001010111110011111111111111111111111111111111111111111111111111111111111111111111111111101011101111000111011111111110010101111,
	240'b101011111111111011011110010111010100111101001110010111101100011101110101010100000101010101010101010101000101000001011000011111111011011111011111111110001111111111111111111111111111111111111110110101000110111001100111111100011111110010101111,
	240'b101011111111111011011101011000101001010010100110101100101111100010110100010110010101010001010101010101010101010101010100010100010101001001100000011101011000111110100011101011001010101110001010010111010100111101101011111100011111110010101111,
	240'b101011111111111011011100011001101110001111110110111010101111110111011000011000000101001101010101010101010101010101010101010101010101010101010011010100010101000001010000010011110100111101010000010100110101001001101011111100011111110010101111,
	240'b101011111111111011011110010110111011111111000101011010111110100110000110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111111011011110010110000111110011101001100001001110101010000011010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111111011011110010111000101010111010000101111001010001101101110010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111111011011110010111000100111010001110111001110110001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101010111100011111110010101111,
	240'b101000011111111011100111011000100101000001011101110111001010000001010000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110010111110001111010110100110,
	240'b100100111111011011111101100110010100111101001101011011000110111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101001110110000111111111110010010010111,
	240'b110000001101001111111111111101011011010010011010100110001001100110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111011111111111011111111111100100010111111,
	240'b111011101100000011100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101100000111110000,
	240'b111110101110111110111110110010111110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110111111101011110001011001001110010001111010111111001,
	240'b111111111111010111100000101000001010000110110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100011001111110110000111110001111111111111110,
	240'b111100101111110011100111101011001010111110110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011010110010101011111001101111010011110011,
	240'b111100001111100011001101110000011101011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111101001010111011110010011110111111110000,
	240'b111100011100011011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001100100011110011,
	240'b110010101100101111111111111111011110010111011000110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011011010110110110001110100111111111111111101100001011001010,
	240'b100101111111001111111111110100111010100110100111101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001011010110110001101001101010110011011110111111111110000110011001,
	240'b100111101111110111110101101100101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001101010111100101101010111010011110111010111111011111001010100100,
	240'b101011101111110011101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001111011011111110110101111101010011010110101111110001111101110101111,
	240'b101011111111110011101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101101011100100111100101110111101010011110110101111110001111101110101111,
	240'b101011111111110011101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110001101111010011000101111101001011010110110011111110001111101110101111,
	240'b101011111111110011101111101011101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111110001011111010010110000111010011101010010110011111110001111101110101111,
	240'b101011111111110011101111101011101010100110101001101010001010011110100111101010001010100010101001101010101010101010101010101010101010101010101010101010101010100110110000111010111111110111101011111110001110101110110110111101111111101110101111,
	240'b101011111111110011101111101011101010011110101101101111111100100111001000110001001011101010110000101010101010011110101001101010101010101010101010101010101010100110101111111001011111110111100010110111101101000010110110111101111111101110101111,
	240'b101011111111110011101111101011001011011111100111111111001111111111111111111111101111101011110011111000011100101010110011101010001010100110101010101010101010101010100111110000001110101110101100101001101010011110110101111110001111101110101111,
	240'b101011111111110011101110101110001110111111111111111111111111111111111111111111111111111111111111111111111111111111110100110101111011010110101000101010011010101010101010101011001011000010101010101010101010100110110101111110001111101110101111,
	240'b101011111111110011101101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011001100101010111010100110101010101010101010100110101010101010101010100110110101111110001111101110101111,
	240'b101011111111101111110011111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111101011000010101000101010101010101010101010101010101010100110110101111110001111101110101111,
	240'b101011111111101111111010111110111111111111111111111111111111111111111111111111111111111111111111111111101111011011110101111110101111111111111111111111111110101010110101101010001010101010101010101010101010100110110101111110001111101110101111,
	240'b101011111111101011111011111110111111111111111111111111111111111111111111111111111111111111111111111111011100100010101111110010011111111011111111111111111111111111101100101101001010100010101010101010101010100110110101111110001111101110101111,
	240'b101011111111101111111001111110101111111111111111111111111111111111111111111111111111111111111111111111111101111110100111101011011110110111111111111111111111111111111111111010001010111110101001101010101010100110110101111110001111101110101111,
	240'b101011111111101111110110111101111111111111111111111111111111111111111111111111111111111111111111111111111111100110111000101001101100110111111111111111111111111111111111111111111101101110101010101010101010100110110101111110001111101110101111,
	240'b101011111111101111110001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111101001111011001011110100111111111111111111111111111111111111110111000101101010001010100110110101111110001111101110101111,
	240'b101011111111110011101110111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101100101010011111010111111111111111111111111111111111111111111111101111101100001010011110110101111110001111101110101111,
	240'b101011111111110011101100110101101111111111111111111111111111111111111111111111111111111111111001110100001100100011101001110011111010011010111000111110011111111111111111111111111111111111111111110100001010011010110101111110001111101110101111,
	240'b101011111111110011101101110001001111110111111111111111111111111111111111111111111111111111110110101100101010010111011011111100001010110110101000111000001111111111111111111111111111111111111111111100011010111110110100111110001111101110101111,
	240'b101011111111110011101110101100111111000011111111111111111111111111111111111111111111111111110110101101001010011111011010111111111100010110100101110000001111110011111111111111111111111111111111111111111100011110110010111110001111101110101111,
	240'b101011111111110011101111101011001101100011111111111111111111111111111111111111111111111111110110101101001010011111011010111111111110010110101010101010111110100011111111111111111111111111111111111111111110001010110100111110001111101110101111,
	240'b101011111111110011101111101011001011101011111010111111111111111111111111111111111111111111111000101101001010011111011011111111111111110110111111101001011100100011111110111111111111111111111111111111111111010110111111111101111111101110101111,
	240'b101011111111110011101111101011101010100111100001111111111111111111111111111111111111010111011111101100011010100011001100111001111110011111001001101001111010111111110001111111111111111111111111111111111111110111001111111101101111101110101111,
	240'b101011111111110011101111101011101010011110111011111110101111111111111111111111111101110010101001101010101010101010101011101010111010101110101011101010101010101011101010111111111111111111111111111111111111111111011111111101011111101110101111,
	240'b101011111111110011101111101011101010100110101001110101101111111111111111111111111101101010100110101010101010101010101001101010001010100010101000101010001010100111101010111111111111111111111111111111111111111111101100111110001111101110101111,
	240'b101011111111110011101111101011101010100110101001101011111110110011111111111111111110111011010001101011111010100011000011110110001101011111010111110101111101011111110101111111111111111111111111111111111111111111110110111110101111101110101111,
	240'b101011111111110011101111101011101010100110101010101010001011101111110110111111111111111111111000101101001010011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110111111101010101111,
	240'b101011111111110011101111101011101010100110101010101010101010100011000011111110001111111111110111101110001010110011011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111101010101111,
	240'b101011111111110011101111101011101010100110101010101010101010101010101000110001001111011111111111111100001110110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111101010101111,
	240'b101011111111110011101111101011101010100110101010101010101010101010101010101010001011111011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111110011111101110101111,
	240'b101011111111110011101111101011101010100110101010101010101010101010101010101010101010100010110011110110111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111101101111101110101111,
	240'b101011111111110011101111101011101010100110101010101010101010110010101011101010101010101010101001101010011100000011100101111111001111111111111111111111111111111111111111111111111111111111111111111111111110101110111011111101111111101110101111,
	240'b101011111111110011101111101011101010011110100110101011111110001110111010101010001010101010101010101010101010100010101100101111111101101111101111111111001111111111111111111111111111111111111110111010011011011110110011111110001111101110101111,
	240'b101011111111110011101111101100001100101011010010110110001111110011011001101011001010100110101010101010101010101010101001101010001010100010101111101110101100011111010001110101011101010111000101101011101010011110110101111110001111101110101111,
	240'b101011111111110011101110101100111111000111111010111101011111111011101100101100001010100110101010101010101010101010101010101010101010101010101001101010001010100010100111101001111010011110101000101010011010100110110101111110001111101110101111,
	240'b101011111111110011101111101011011101111111100010101101011111010011000011101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110001111101110101111,
	240'b101011111111110011101111101011001011111011110100110000101111010111000001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110001111101110101111,
	240'b101011111111110011101111101011011010101011100111110111011101000110110111101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110001111101110101111,
	240'b101011111111110011101111101011101010011111000111111100111011000110101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110110101111110001111101110101111,
	240'b101000011111110111110100101100001010100010101110111011101100111110101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010111000111111001111010010100110,
	240'b100100111111011011111110110011001010011110100110101101101011011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010100111010111111111111110010010010111,
	240'b110000001101001111111111111110101101101011001101110011001100110011001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011101111111111101111111111100100010111111,
	240'b111011101100000011100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101100000111110000,
	240'b111110101110111110111110110010111110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101011110001011001001110010001111010111111001,
	240'b111111111111010111100000101000001010000110110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100011001111110110000111110001111111111111110,
	240'b111100101111110011100111101011001010111110110110101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101011010110010101011111001101111010011110011,
	240'b111100001111100011001101110000011101011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111101001010111011110010011110111111110000,
	240'b111100011100011011011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001100100011110011,
	240'b110010101100101111111111111110111100101010110001101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001010111010101110101100101101001111111111111111101100001011001010,
	240'b100101111111001111111110101010000101010001010000010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010110101101100010010011100101101010111110111111111110001010011001,
	240'b100111101111111011101011011001010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100011010110011001011010101100100111101110110111110101111001110100100,
	240'b101011101111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000111000011101101011111010100111001101010111100011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011011011001001001111001010101111100100111101101010111100011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100011011110100110001011111010010110101101100111111100011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100011001110100001100001110100111010100101100110111100011111110010101111,
	240'b101011111111111011011110010111010101010001010100010100010100111101001111010100000101000101010011010101000101010101010101010101010101010101010101010101010101001101100001110101111111101011010110111100011101100001101110111100001111110010101111,
	240'b101011111111111011011110010111010101000001011011100000001001010010010001100010000111011001100010010101010101000001010011010101010101010101010101010101010101001101011110110011001111101011000100101111101010000101101110111100001111110010101111,
	240'b101011111111111011011110010110010111000011001110111110011111111111111111111111011111010011100111110000111001011001100111010100100101001001010101010101010101010101010000100000101101011001011000010011100100111001101011111100011111110010101111,
	240'b101011111111111011011011011100011101111111111111111111111111111111111111111111111111111111111111111111111111111111101000101011110110101001010001010101000101010101010101010110010110000101010110010101010101001001101011111100011111110010101111,
	240'b101011111111111011011011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010011001010101110101001001010101010101000101001101010101010101010101001001101011111100011111110010101111,
	240'b101011111111110011100111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111100110001101010001010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111101111110100111101101111111111111111111111111111111111111111111111111111111111111111111111011110110111101011111101101111111111111111111111111101010101101010010100010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111101111110101111101111111111111111111111111111111111111111111111111111111111111111111111110111001000001011111100101001111110111111111111111111111111111011001011010010101000101010101010101010101001001101011111100011111110010101111,
	240'b101011111111101111110010111101001111111111111111111111111111111111111111111111111111111111111111111111111011111001001111010110111101101111111111111111111111111111111111110100000101111101010011010101010101001001101011111100011111110010101111,
	240'b101011111111110011101100111100001111111111111111111111111111111111111111111111111111111111111111111111111111001101110001010011001001110011111111111111111111111111111111111111111011011001010100010101000101001001101011111100011111110010101111,
	240'b101011111111110111100011111001101111111111111111111111111111111111111111111111111111111111111111111111111111111110101110010011100110010111101000111111111111111111111111111111111111101010001011010100000101001001101011111100011111110010101111,
	240'b101011111111110111011101110100001111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011001010100111010101110111111111111111111111111111111111111111111011111011000010101000001101011111100011111110010101111,
	240'b101011111111111011011001101011101111111111111111111111111111111111111111111111111111111111110100101000101001000111010011100111110100110001110010111100111111111111111111111111111111111111111111101000100100110101101011111100011111110010101111,
	240'b101011111111111011011001100010011111101111111111111111111111111111111111111111111111111111101110011001100100101010110110111000000101110001010010110000001111111111111111111111111111111111111111111000110101111101101000111100011111110010101111,
	240'b101011111111111011011100011001111110000111111111111111111111111111111111111111111111111111101110011010100100111110110101111111111000101101001011100000001111101011111111111111111111111111111111111111101000111101100110111100011111110010101111,
	240'b101011111111111011011110010110011011000011111111111111111111111111111111111111111111111111101110011010100100111110110100111111111100101101010101010101111101000111111111111111111111111111111111111111111100010101101010111100001111110010101111,
	240'b101011111111111011011110010110010111010111110110111111111111111111111111111111111111111111110010011010110100111110110111111111111111110001111110010011001001000111111101111111111111111111111111111111111110101101111111111011101111110010101111,
	240'b101011111111111011011110010111000101001111000010111111111111111111111111111111111110101111000000011001000101000110011000110100001101000110010100010100000110000011100100111111111111111111111111111111111111110010011110111011001111110010101111,
	240'b101011111111111011011110010111010100111101110111111101011111111111111111111111111011011101010011010101010101010101010111010110000101100001011000010101000101011011010100111111111111111111111111111111111111111111000000111011001111110010101111,
	240'b101011111111111011011110010111010101001101010010101011011111111111111111111111111011010001001100010101000101010101010011010100010101000101010001010100010101010011010100111111111111111111111111111111111111111111011001111100001111110010101111,
	240'b101011111111111011011110010111010101010001010011010111111101100011111111111111111101111010100100011000000101001010001000101100011011000010110000101011111011000011101011111111111111111111111111111111111111111111101101111101001111101110101111,
	240'b101011111111111011011110010111010101010001010101010100010111011011101100111111111111111111110010011010010100110110110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101111111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101000010000110111100011111111111101111011100100101100010111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110001111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010001100010101110111011111111111000011101101111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111110001111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101010101010101010100000111110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111101001111101110101111,
	240'b101011111111111011011110010111010101010001010101010101010101010001010101010101010101000101100111101110001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111000111011011111110010101111,
	240'b101011111111111011011110010111010101010001010101010101010101100101010110010101010101010101010010010101001000000111001010111110011111111111111111111111111111111111111111111111111111111111111111111111111101011101111000111011111111110010101111,
	240'b101011111111111011011110010111010100111101001110010111101100011101110101010100000101010101010101010101000101000001011000011111111011011111011111111110001111111111111111111111111111111111111110110101000110111001100111111100011111110010101111,
	240'b101011111111111011011101011000101001010010100110101100101111100010110100010110010101010001010101010101010101010101010100010100010101001001100000011101011000111110100011101011001010101110001010010111010100111101101011111100011111110010101111,
	240'b101011111111111011011100011001101110001111110110111010101111110111011000011000000101001101010101010101010101010101010101010101010101010101010011010100010101000001010000010011110100111101010000010100110101001001101011111100011111110010101111,
	240'b101011111111111011011110010110111011111111000101011010111110100110000110010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111111011011110010110000111110011101001100001001110101010000011010100000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111111011011110010111000101010111010000101111001010001101101110010100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101011111100011111110010101111,
	240'b101011111111111011011110010111000100111010001110111001110110001101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001101010111100011111110010101111,
	240'b101000011111111011100111011000100101000001011101110111001010000001010000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101110010111110001111010110100110,
	240'b100100111111011011111101100110010100111101001101011011000110111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110100111101001111010011110101001110110000111111111110010010010111,
	240'b110000001101001111111111111101011011010010011010100110001001100110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111011111111111011111111111100100010111111,
	240'b111011101100000011100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101101100000111110000,
	240'b111110101110111110111110110010111110011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110111111101011110001011001001110010001111010111111001,
	240'b111111111111010111100000101000001010000110110011101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101100011001111110110000111110001111111111111110,
};
assign data = picture[addr];
endmodule