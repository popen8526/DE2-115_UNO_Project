module blue_nine(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111111111111110111011101100110011010000110111001101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110001001110110100110111100111111111111111111,
	240'b111111111110110010110111110101001110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011010000110000011111011011111111,
	240'b111110001011111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100001111111100,
	240'b110010011101110011111111111011101010110110010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001000110001111100100111011010011110100111111111101010011001011,
	240'b101000001111101111111001100010100100111001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011100110100110000101011001010100110110011010111111101111011110010111,
	240'b101100101111111111011101010110010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100001011110110011110101111010000111100101100001111010101111111010100111,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110110001100011101110111110100011100110001100000111000001111111110110110,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010101000110001000010100110101110000101101000110111111111111110110110,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111011001101001010001100110111101100001001011110111000011111111110110110,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010001111000011110000110101100110110101011100111000011111111110110110,
	240'b110000101111111111010010010101100101010001010011010100000101000101010000010011110101000001010010010101000101010101010101010101010101010101010101010101010101001101100011111001101010001101101101011100110101100101011110111000011111111110110110,
	240'b110000101111111111010010010101100101000001100101100100001010010110100011100110001000010101101110010110010101000101010001010101000101010101010101010101010101010101010100101110111110110010110111111010001001001001011011111000011111111110110111,
	240'b110000101111111111010010010100111000010111100001111111111111111111111111111111111111110011110000110101001010100101110110010101010101000101010101010101010101010101010011011000111011100011011101101100100110000001011101111000011111111110110111,
	240'b110000101111111111001110011110111111000011111111111111111111111111111111111111111111111111111111111111111111111111110100110000100111100101010010010100110101010101010101010100110101010001011011010100110101000101011111111000011111111110110111,
	240'b110000101111111111010011110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110101100010111100101000101010101010101010101010001010100010101010101001101011111111000011111111110110111,
	240'b110000101111111111101001111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000110111001010001010101010101010101010101010101010101001101011111111000011111111110110111,
	240'b110000101111111111110100111111011111111111111111111111111111111111111111111111111111111111111111111111111111100011101010111010111111101011111111111111111110001101111001010100000101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111110100111111011111111111111111111111111111111111111111111111111111111111111101110000110111110001100001011000111000001111001101111111111111111111101000011110000101000101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111110011111111011111111111111111111111111111111111111111111111111111111010101110010101100100111101001101010011100100111001011011101111101111111111111111111000010110101001010001010101010101001101011111111000011111111110110110,
	240'b110000101111111111101100111101011111111111111111111111111111111111111111111111111101011001011011010100000110000110001101100010010101110001001111011001001110001111111111111111111100101001011010010101000101001101011111111000011111111110110110,
	240'b110000101111111111100001111010001111111111111111111111111111111111111111111111111001100001001101011000001100110111111111111111101011111101011010010011101010101011111111111111111111111110100000010100010101001101011111111000011111111110110110,
	240'b110000101111111111010100110101011111111111111111111111111111111111111111111110010111011101001100100101001111111111111111111111111111111010000010010010111000100011111110111111111111111111101101011011100101000001011111111000011111111110110111,
	240'b110000101111111111001110101101001111111111111111111111111111111111111111111101010110110101001100101001111111111111111111111111111111111110010010010010111000000111111100111111111111111111111111101101110101000101011110111000011111111110110111,
	240'b110000101111111111001101100011011111111011111111111111111111111111111111111101010110110001001110100000111111110011111111111111111111010101110011010011001001000011111111111111111111111111111111111100010110110101011011111000011111111110110111,
	240'b110000101111111111001111011001111110101011111111111111111111111111111111111101010110110001010001010101101010010111101010111001101001011101010011010100011011110011111111111111111111111111111111111111111010011001011010111000011111111110110111,
	240'b110000101111111111010001010101001011110011111111111111111111111111111111111101010110110001010010010100110101010001100100011000100101001101001110011110111111001111111111111111111111111111111111111111111101100101100101111000001111111110110111,
	240'b110000101111111111010010010100100111111011111010111111111111111111111111111101010110110001010010010110000101001001001101010011010101000001111000111000011111111111111111111111111111111111111111111111111111011110000011110111011111111110110111,
	240'b110000101111111111010010010101010101011111001011111111111111111111111111111101010110110001001110100101111010111110001001100011001011001111110000111111111111111111111111111111111111111111111111111111111111111110100111110111001111111110110110,
	240'b110000101111111111010010010101100101000001111110111110001111111111111111111110000111011001001100100110101111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111001001110111111111111010110110,
	240'b110000101111111111010010010101100101001101010100101101011111111111111111111111101001010001001101011001001101011111111111111111111100001110000010110010101111101011111111111111111111111111111111111111111111111111100011111001001111111010110110,
	240'b110000101111111111010010010101100101010001010010011001001101111111111111111111111101001001011001010100000110011110011010100100110101111101001100011001101110100111111111111111111111111111111111111111111111111111101110111011001111110110110110,
	240'b110000101111111111010010010101100101010001010101010100010111110011110000111111111111110110100101010100110100111101001111010011110100111101010111101101001111111011111111111111111111111111111111111111111111111111110011111100101111110110110110,
	240'b110000101111111111010010010101100101010001010101010101010101000010001101111101001111111111111011101110010111011001100011011000110111101011000011111111101111111111111111111111111111111111111111111111111111111111110110111101011111110010110111,
	240'b110000101111111111010010010101100101010001010101010101010101010101010001100100001111001011111111111000111011010010100010101000101011011111101011111111111111111111111111111111111111111111111111111111111111111111110110111101011111110010110111,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010100011000000111100110110001000111111010000010100000100111111011001110111111111111111111111111111111111111111111111111111111111111111111101101111010111111110110110111,
	240'b110000101111111111010010010101100101010001010101010101000101010101010101010101010101000001101100110000011111101011111111111111101111110111111110111111111111111111111111111111111111111111111111111111111111111111000100110111101111111110110111,
	240'b110000101111111111010010010101100101001001010010010101110101001001010100010101010101010101010010010101111000101011010011111110111111111111111111111111111111111111111111111111111111111111111111111111111110100101111010110111101111111110110111,
	240'b110000101111111111010010010101010110001010101110110011111010001001011010010101000101010101010101010101000101000001011010100000111011101111100100111110001111111111111111111111111111111111111111111000111000000001011011111000011111111110110110,
	240'b110000101111111111010010010100111010001111101101110001111111010010100001010100010101010101010101010101010101010101010100010100010101001101100010011111011001010010101000101100111011001110011000011010000101000001011111111000011111111110110110,
	240'b110000101111111111010010010101010110001101110110011000111011010111011100010101110101010001010101010101010101010101010101010101010101010001010011010100010101000001010001010100100101001001010000010100100101001101011111111000011111111110110110,
	240'b110000101111111111010010010100110111001011010101111011011110110011100000010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111010001010110011101000011011001100110111110011011100001010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111001111011001111110111110000101010000101010001011100100010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111010000010111101110001010110111011010111100111011001101010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110111,
	240'b101101001111111111011011010101011001001011110011111100111110110001111111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100011111010001111111110101001,
	240'b100111111111110011110111100000100100110101110101100100010110110001001110010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111010010011111111011111100010010110,
	240'b110001011110000111111111111010011001111110000101100001001000011010001001100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010011010011111110000111111111101011111000101,
	240'b111101101011111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011100001011111011,
	240'b111101101110010010111110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011011000101110101110100011110110,
	240'b111011101111011111101101100110101001000110101011101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010101000110110011100111001001111000111101110,
	240'b111111111111110111011101100110011010000110111001101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110001001110110100110111100111111111111111111,
	240'b111111111110110010110111110101001110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011010000110000011111011011111111,
	240'b111110001011111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100001111111100,
	240'b110010011101110011111111111011101010110110010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001000110001111100100111011010011110100111111111101010011001011,
	240'b101000001111101111111001100010100100111001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010011100110100110000101011001010100110110011010111111101111011110010111,
	240'b101100101111111111011101010110010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100001011110110011110101111010000111100101100001111010101111111010100111,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011010110110001100011101110111110100011100110001100000111000001111111110110110,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010101000110001000010100110101110000101101000110111111111111110110110,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111011001101001010001100110111101100001001011110111000011111111110110110,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100111111010001111000011110000110101100110110101011100111000011111111110110110,
	240'b110000101111111111010010010101100101010001010011010100000101000101010000010011110101000001010010010101000101010101010101010101010101010101010101010101010101001101100011111001101010001101101101011100110101100101011110111000011111111110110110,
	240'b110000101111111111010010010101100101000001100101100100001010010110100011100110001000010101101110010110010101000101010001010101000101010101010101010101010101010101010100101110111110110010110111111010001001001001011011111000011111111110110111,
	240'b110000101111111111010010010100111000010111100001111111111111111111111111111111111111110011110000110101001010100101110110010101010101000101010101010101010101010101010011011000111011100011011101101100100110000001011101111000011111111110110111,
	240'b110000101111111111001110011110111111000011111111111111111111111111111111111111111111111111111111111111111111111111110100110000100111100101010010010100110101010101010101010100110101010001011011010100110101000101011111111000011111111110110111,
	240'b110000101111111111010011110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110101100010111100101000101010101010101010101010001010100010101010101001101011111111000011111111110110111,
	240'b110000101111111111101001111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000110111001010001010101010101010101010101010101010101001101011111111000011111111110110111,
	240'b110000101111111111110100111111011111111111111111111111111111111111111111111111111111111111111111111111111111100011101010111010111111101011111111111111111110001101111001010100000101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111110100111111011111111111111111111111111111111111111111111111111111111111111101110000110111110001100001011000111000001111001101111111111111111111101000011110000101000101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111110011111111011111111111111111111111111111111111111111111111111111111010101110010101100100111101001101010011100100111001011011101111101111111111111111111000010110101001010001010101010101001101011111111000011111111110110110,
	240'b110000101111111111101100111101011111111111111111111111111111111111111111111111111101011001011011010100000110000110001101100010010101110001001111011001001110001111111111111111111100101001011010010101000101001101011111111000011111111110110110,
	240'b110000101111111111100001111010001111111111111111111111111111111111111111111111111001100001001101011000001100110111111111111111101011111101011010010011101010101011111111111111111111111110100000010100010101001101011111111000011111111110110110,
	240'b110000101111111111010100110101011111111111111111111111111111111111111111111110010111011101001100100101001111111111111111111111111111111010000010010010111000100011111110111111111111111111101101011011100101000001011111111000011111111110110111,
	240'b110000101111111111001110101101001111111111111111111111111111111111111111111101010110110101001100101001111111111111111111111111111111111110010010010010111000000111111100111111111111111111111111101101110101000101011110111000011111111110110111,
	240'b110000101111111111001101100011011111111011111111111111111111111111111111111101010110110001001110100000111111110011111111111111111111010101110011010011001001000011111111111111111111111111111111111100010110110101011011111000011111111110110111,
	240'b110000101111111111001111011001111110101011111111111111111111111111111111111101010110110001010001010101101010010111101010111001101001011101010011010100011011110011111111111111111111111111111111111111111010011001011010111000011111111110110111,
	240'b110000101111111111010001010101001011110011111111111111111111111111111111111101010110110001010010010100110101010001100100011000100101001101001110011110111111001111111111111111111111111111111111111111111101100101100101111000001111111110110111,
	240'b110000101111111111010010010100100111111011111010111111111111111111111111111101010110110001010010010110000101001001001101010011010101000001111000111000011111111111111111111111111111111111111111111111111111011110000011110111011111111110110111,
	240'b110000101111111111010010010101010101011111001011111111111111111111111111111101010110110001001110100101111010111110001001100011001011001111110000111111111111111111111111111111111111111111111111111111111111111110100111110111001111111110110110,
	240'b110000101111111111010010010101100101000001111110111110001111111111111111111110000111011001001100100110101111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111001001110111111111111010110110,
	240'b110000101111111111010010010101100101001101010100101101011111111111111111111111101001010001001101011001001101011111111111111111111100001110000010110010101111101011111111111111111111111111111111111111111111111111100011111001001111111010110110,
	240'b110000101111111111010010010101100101010001010010011001001101111111111111111111111101001001011001010100000110011110011010100100110101111101001100011001101110100111111111111111111111111111111111111111111111111111101110111011001111110110110110,
	240'b110000101111111111010010010101100101010001010101010100010111110011110000111111111111110110100101010100110100111101001111010011110100111101010111101101001111111011111111111111111111111111111111111111111111111111110011111100101111110110110110,
	240'b110000101111111111010010010101100101010001010101010101010101000010001101111101001111111111111011101110010111011001100011011000110111101011000011111111101111111111111111111111111111111111111111111111111111111111110110111101011111110010110111,
	240'b110000101111111111010010010101100101010001010101010101010101010101010001100100001111001011111111111000111011010010100010101000101011011111101011111111111111111111111111111111111111111111111111111111111111111111110110111101011111110010110111,
	240'b110000101111111111010010010101100101010001010101010101010101010101010101010100011000000111100110110001000111111010000010100000100111111011001110111111111111111111111111111111111111111111111111111111111111111111101101111010111111110110110111,
	240'b110000101111111111010010010101100101010001010101010101000101010101010101010101010101000001101100110000011111101011111111111111101111110111111110111111111111111111111111111111111111111111111111111111111111111111000100110111101111111110110111,
	240'b110000101111111111010010010101100101001001010010010101110101001001010100010101010101010101010010010101111000101011010011111110111111111111111111111111111111111111111111111111111111111111111111111111111110100101111010110111101111111110110111,
	240'b110000101111111111010010010101010110001010101110110011111010001001011010010101000101010101010101010101000101000001011010100000111011101111100100111110001111111111111111111111111111111111111111111000111000000001011011111000011111111110110110,
	240'b110000101111111111010010010100111010001111101101110001111111010010100001010100010101010101010101010101010101010101010100010100010101001101100010011111011001010010101000101100111011001110011000011010000101000001011111111000011111111110110110,
	240'b110000101111111111010010010101010110001101110110011000111011010111011100010101110101010001010101010101010101010101010101010101010101010001010011010100010101000001010001010100100101001001010000010100100101001101011111111000011111111110110110,
	240'b110000101111111111010010010100110111001011010101111011011110110011100000010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111010001010110011101000011011001100110111110011011100001010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111001111011001111110111110000101010000101010001011100100010110010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110110,
	240'b110000101111111111010000010111101110001010110111011010111100111011001101010101000101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011111111000011111111110110111,
	240'b101101001111111111011011010101011001001011110011111100111110110001111111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100011111010001111111110101001,
	240'b100111111111110011110111100000100100110101110101100100010110110001001110010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000100111010010011111111011111100010010110,
	240'b110001011110000111111111111010011001111110000101100001001000011010001001100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010011010011111110000111111111101011111000101,
	240'b111101101011111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011100001011111011,
	240'b111101101110010010111110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011011000101110101110100011110110,
	240'b111011101111011111101101100110101001000110101011101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010101000110110011100111001001111000111101110,
	240'b111111111111110111011101100110011010000110111001101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110101011101010111010101110001001110110100110111100111111111111111111,
	240'b111111111110110010110111110101001110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110110011010000110000011111011011111111,
	240'b111110001011111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100001111111100,
	240'b110010011101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010011001011,
	240'b101000001111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010010111,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010100111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110110,
	240'b110000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111,
	240'b101101001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010101001,
	240'b100111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110010110,
	240'b110001011110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111000101,
	240'b111101101011111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010011100001011111011,
	240'b111101101110010010111110110111101110111011101110111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101110111011011000101110101110100011110110,
	240'b111011101111011111101101100110101001000110101011101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010101000110110011100111001001111000111101110,
};
assign data = picture[addr];
endmodule