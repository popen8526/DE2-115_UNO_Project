// audio.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module audio (
		output wire  altpll_0_c0_clk,                      //                    altpll_0_c0.clk
		input  wire  altpll_0_inclk_interface_clk,         //       altpll_0_inclk_interface.clk
		input  wire  altpll_0_inclk_interface_reset_reset, // altpll_0_inclk_interface_reset.reset
		output wire  altpll_1_c0_clk,                      //                    altpll_1_c0.clk
		input  wire  altpll_1_inclk_interface_clk,         //       altpll_1_inclk_interface.clk
		input  wire  altpll_1_inclk_interface_reset_reset  // altpll_1_inclk_interface_reset.reset
	);

	audio_altpll_0 altpll_0 (
		.clk       (altpll_0_inclk_interface_clk),         //       inclk_interface.clk
		.reset     (altpll_0_inclk_interface_reset_reset), // inclk_interface_reset.reset
		.read      (),                                     //             pll_slave.read
		.write     (),                                     //                      .write
		.address   (),                                     //                      .address
		.readdata  (),                                     //                      .readdata
		.writedata (),                                     //                      .writedata
		.c0        (altpll_0_c0_clk),                      //                    c0.clk
		.areset    (),                                     //        areset_conduit.export
		.locked    (),                                     //        locked_conduit.export
		.phasedone ()                                      //     phasedone_conduit.export
	);

	audio_altpll_1 altpll_1 (
		.clk       (altpll_1_inclk_interface_clk),         //       inclk_interface.clk
		.reset     (altpll_1_inclk_interface_reset_reset), // inclk_interface_reset.reset
		.read      (),                                     //             pll_slave.read
		.write     (),                                     //                      .write
		.address   (),                                     //                      .address
		.readdata  (),                                     //                      .readdata
		.writedata (),                                     //                      .writedata
		.c0        (altpll_1_c0_clk),                      //                    c0.clk
		.areset    (),                                     //        areset_conduit.export
		.locked    (),                                     //        locked_conduit.export
		.phasedone ()                                      //     phasedone_conduit.export
	);

endmodule
