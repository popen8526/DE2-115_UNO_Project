module wild(
	input [7:0] addr,
	output [239:0] data
);
parameter [0:149][239:0] picture = {
	240'b111010011111110111001001011110001001001110101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010001000010010001101111010011111110111111010,
	240'b111100001111000010111010110011011110001111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010111101110111000110110010101111110011111111,
	240'b111001001100000011101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100101111111111,
	240'b101110101110001011111111111001101000101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111001101010011010010110100101101110011100011010011011111010111111111100101111001111,
	240'b101011101111110111110001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001111011001100011010000000000000000000000001110001001111111111110101010011110,
	240'b101100001111111110111000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011010010000110000001111100010100010000110000000000000101000111100001111101110101010,
	240'b101100001111111110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111101100111011010111111001011111111101100100000101100011001111000101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101001110111010010011010101011111000111110100110000100010101111000101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110101110111000011100010110011010100111101111011001100100000111000011111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101101100001110010000000001111000111111111101111000110101110111101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011011110010100111000101000111000001110001100110100110111111111111110110001,
	240'b101100011111111110100010000000000000001101000001011110011000110110011111100100100111010101000011000110100000000000000000000000000000000000000000000000000000000000000000000011000101011101110101101010110110101000011011111000101111111110110001,
	240'b101100011111111110100000000010100111011010010111011011110111011011110001111111111111111111111011110111011010000101001100000010110000000000000000000000000000000000000000000000000000000000000111000010010000000000011011111000101111111110110001,
	240'b101100011111111110100000011010111000100001010010010100100100111110100010111111111111111111111111111111111111111111111100110000000100111100000010000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111000110100101000101010001010100010101010101001101100010111000011111111111111111111111111111111111111111111111111111100010100001001000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111100111011101000101000101010101010101010101010101010000100101101111111011111111111111111111111111111111111111111111111111111111110101000100000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111101001011000010101001101010101010101010101010101010011010111011101100011111111111111111111111111111111111111111111111111111111111111111110100101001111000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111100111010111110101001101010101010101010101010101010101010100001000110011111100111111111111111111111111111111111111111111111111111111111111111111101101010011110000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111101010011001000101001101010101010101010101010101010101010101000101100011001110111111111111111111111111111111111111111111111111111111111111111111111111111001100011010000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111101001011010110101001001010101010101010101010101010101010101010101000010000010111110011111111111111111111111111111111111111111111111111111111111111111111111111100010100010011000000000000000000011100111000101111111110110001,
	240'b101100001111111111100001011101110101000101010101010101010101010101010101010101010101010001010101110001001111111111111111111111111111111111111111111111111111111111111111111111111111111110001010000000000000000000011100111000101111111110110001,
	240'b101100001111111111010100100001110101000101010101010101010101010101010101010101010101010101010001011110001111010111111111111111111111111111111111111111111111111111111111111111111111111111110001001110000000000000011100111000101111111110110001,
	240'b101100011111111110111100100011110101010001010101010101010101010101010101010101010101010101010101010100101011100111111111111111111111111111111111111111111111111111111111111111111111111111111111101010100000000100011011111000101111111110110001,
	240'b101100011111111110100101100001000110000101010100010101010101010101010101010101010101010101010101010100010110111111110000111111111111111111111111111111111111111111111111111111111111111111111111111101010011010000010101111000101111111110110001,
	240'b101100011111111110011100010110110111111001011000010110110101101101011011010110110101101101011011010110110101011110110010111111111111111111111111111111111111111111111111111111111111111111111111111111111001000000010111111000101111111110110001,
	240'b101100011111111110011110001001110111101000011011000111010001110100011101000111010001110100011101000111010001101100110011110111101111111111111111111111111111111111111111111111111111111111111111111111111101011100110001110111111111111110110001,
	240'b101100011111111110100010000000110111000100010111000000000000000000000000000000000000000000000000000000000000000000000000011101001111111111111111111111111111111111111111111111111111111111111111111111111111100101100111110110111111111110110001,
	240'b101100011111111110100010000000000011111001011101000000000000000000000000000000000000000000000000000000000000000000000000000101001101001011111111111111111111111111111111111111111111111111111111111111111111111110100011110110111111111110110001,
	240'b101100001111111110100010000000000000011001110111000111100000000000000000000000000000000000000000000000000000000000000000000000000110010011111110111111111111111111111111111111111111111111111111111111111111111111010111111001011111111010110001,
	240'b101100001111111110100010000000000000000000110010011011110000001000000000000000000000000000000000000000000000000000000000000000000000110111000101111111111111111111111111111111111111111111111111111111111111111111110011111011011111110110110001,
	240'b101100001111111110100010000000000000000000000000011001000100100000000000000000000000000000000000000000000000000000000000000000000000000001010011111110111111111111111111111111111111111111111111111111111111111111110111111101001111110010110001,
	240'b101100001111111110100010000000000000000000000000000011000111101000101011000000000000000000000000000000000000000000000000000000000000000000000111101101111111111111111111111111111111111111111111111111111111111111111100111110111111110010110001,
	240'b101100001111111110100010000000000000000000000000000000000001110101111111001000010000000000000000000000000000000000000000000000000000000000000000010001001111011111111111111111111111111111111111111111111111111111111110111111011111110010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000100111100000010010100000000000000000000000000000000000000000000000000000000000000001001010100011111111111111111111111111111111111111111111111111111110111111101111110010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000001001001000001000111111000000000000000000000000000000000000000000000000000000000011011011110001111111111111111111111111111111111111111111111011111110001111110010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000001001101110001011010000001010000000000000000000000000000000000000000000000000110011000111111111111111111111111111111111111111111100010111010011111111010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000000000000000010010001011000000001010101000101100000000000000000000000000000000000101001111010011111111111111111111111111111101101111100110111001111111110110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010010011111100110101100111101000111000000100000000000100001111111111111111111111111001000100000011111111000011111111110110001,
	240'b101100001111111110100001000000110101000001110111010100010000110100000000000000000000000000000000000000000000000000000000000010100011001101011110011101100111101001110011100010011110000010111110010111100000001100011010111000101111111110110001,
	240'b101100001111111110011100001111001001010010101000111111101100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100011111001000100001110100001001000000000000000000011100111000101111111110110001,
	240'b101100001111111110011011010100100111101001011001110111011111111111010011001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111110011100001110111000010101001000100010101111011111111110100011110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111110100000000100110111110000010100000101101011101111111101110110110001011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111110100001000000000101001001010110000000000100101011111010111110100011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111000101111111110110001,
	240'b101100011111111110101011000000000000011001101010011001010010000110111100111111010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010011111111010101110,
	240'b101011101111111111100000000111110000000000000000001111100110110110010111011110010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100111111011111000010011110,
	240'b101100001110111011111111101110010100010000101110001010110011000100110101001011010010111100110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000101111111100010111111111101010110110111,
	240'b110101101100010011111100111111111111100011101101111011011110110111101100111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101111111111111111111011011100000111110111,
	240'b111011101101101111000001111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100000101111001110110111111110,
	240'b111000001111011011011101101001101010001110101010101010111010101010101010101010101010101010101010101010111010101110101011101010111010101010101010101010101010101010101010101010101010101110101011101010011010000110101101111001101111010011110001,
	240'b111010011111110111001001011110001001001110101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010001000010010001101111010011111110111111010,
	240'b111100001111000010111010110011011110001111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010111101110111000110110010101111110011111111,
	240'b111001001100000011101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100101111111111,
	240'b101110101110001011111111111001101000101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111001101010011010100110101001101110011100011010011011111010111111111100101111001111,
	240'b101011101111110111110001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001110010111110011010100000000000000000000001110001001111111111110101010011110,
	240'b101100001111111110111000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011110010010011101001001001110000110000110110000000000101000111100001111101110101010,
	240'b101100001111111110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111101101010010010100100111101110110100011100000110100011001111000101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101001111000010011010100110001001100100000000101101000010110111000101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100110101011100011001000011110000101100101011001100100100011111000011111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001110001101010101010100000101011011011010000110111110111101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100100111100011110101110101011001011100100110110110111111111111110110001,
	240'b101100011111111110100010000000000000001101000001011110011000011110000100011110110110100101000101000111100000000100000000000000000000000000000000000000000000000000000000000010010101101110011101101100000110000100011011111000101111111110110001,
	240'b101100011111111110100000000010100111011010010111011100010110100101101101011011100111101010001101100110001000010101001100000011110000000000000000000000000000000000000000000000000000000000000011000010010000000000011011111000101111111110110001,
	240'b101100011111111110100000011010111000100001010010010100100101010001011111010101000101001001010001010101100110101010001110100101100100111100000110000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111000110100101000101010001010100010101010101010001011011010111010101010001010101010101010101001101010001011000101001000110001001001001010000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111100111011101000101000101010101010101010101010101010101011000000101011101010101010101010101010101010101010100110101001001110100100111010100001000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111101001011000010101001101010101010101010101010101010100010110100101111001010100010101010101010101010101010101010101010101010001011000011001101001001111000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111100111010111110101001101010101010101010101010101010101010101010110000001011000010101010101010101010101010101010101010101010101010100110101101010011001010011110000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111101010011001000101001101010101010101010101010101010101010101010101100001011111010101010101010101010101010101010101010101010101010101010101001101011011100111010011100000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111101001011010110101001001010101010101010101010101010101010101010101010001011111010110010101010001010101010101010101010101010101010101010101010101010010011001001001010100010111000000000000000000011100111000101111111110110001,
	240'b101100001111111111100001011101110101000101010101010101010101010101010101010101010101010101010111011000000101010101010101010101010101010101010101010101010101010101010101010100010111101001111001000000100000000000011100111000101111111110110001,
	240'b101100001111111111010100100001110101000101010101010101010101010101010101010101010101010101010100010111100101101001010101010101010101010101010101010101010101010101010101010101010101001110010100001110100000000000011100111000101111111110110001,
	240'b101100011111111110111100100011110101010001010101010101010101010101010101010101010101010101010101010101110110000001010101010101010101010101010101010101010101010101010101010101010101001101100111100010010000010000011011111000101111111110110001,
	240'b101100011111111110100101100001000110000001010011010101000101010001010100010101000101010001010100010100110101110001011010010100110101010001010100010101000101010001010100010101000101010001010001100011100011011000010110111000101111111110110001,
	240'b101100011111111110011100010110111000000001011000010110110101101101011011010110110101101101011011010110110101110101100110010111000101101101011011010110110101101101011011010110110101101101011001011100100111100000011010111000101111111110110001,
	240'b101100011111111110011110001000111011001110011100100110111001101110011011100110111001101110011011100110111001101110011111100111111001101110011011100110111001101110011011100110111001101110011011100111101010111000110100110111111111111110110001,
	240'b101100011111111110100010000000011001000110111010101010111010110010101100101011001010110010101100101011001010110010101100101100101010110110101100101011001010110010101100101011001010110010101100101010111011111001100110110110111111111110110001,
	240'b101100011111111110100010000000000011110011000011101010101010101010101010101010101010101010101010101010101010101010101010101011011010111010101010101010101010101010101010101010101010101010101010101010011011011010011000110111011111111110110001,
	240'b101100001111111110100010000000000000010010010100101110101010100110101010101010101010101010101010101010101010101010101010101010101011000010101011101010101010101010101010101010101010101010101010101010101010111010111110111001111111111010110001,
	240'b101100001111111110100010000000000000000000101110110000001010110110101010101010101010101010101010101010101010101010101010101010101010110010101111101010101010101010101010101010101010101010101010101010101010100111001101111100001111110110110001,
	240'b101100001111111110100010000000000000000000000000011011001100010010101001101010101010101010101010101010101010101010101010101010101010101010101111101010111010101010101010101010101010101010101010101010101010100011000111111101101111110110110001,
	240'b101100001111111110100010000000000000000000000000000010011001010110111110101010001010101010101010101010101010101010101010101010101010101010101100101011111010101010101010101010101010101010101010101010101010100011000011111110101111110010110001,
	240'b101100001111111110100010000000000000000000000000000000000001100110101010101110101010100010101010101010101010101010101010101010101010101010101010101011111010110010101010101010101010101010101010101010101010100011000010111111001111110010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000100011101011101011110110101000101010101010101010101010101010101010101010101010101010111010111110101010101010101010101010101010101010101010100011000001111111011111110010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000111111010001111000010101010111010100110101010101010101010101010101010101010101010111110101100101010101010101010101010101010101010100011001000111110001111110010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000001000001111111110001101011010110101001101010011010101010101010101010101010101110110000101010101010101010101010101010011010110111000110111010111111111010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000000000000000000010001001010100011000110101101101010101010101001101010011010101010101110101011011010101010101001101010101100001101111001110111001111111110110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001010100101000011100001111000001101110011011000110101110101100011010110010110011110001110111111100100000111000011111111110110001,
	240'b101100001111111110100001000000110101000001110000010011100001000100000000000000000000000000000000000000000000000000000000000001100011000001100101100100101010100110111010110000111100000010101000010110110000010000011001111000101111111110110001,
	240'b101100001111111110011100001111001001100001101110100010111001010100110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100011010001000010001111100001011000000000000000000011100111000101111111110110001,
	240'b101100001111111110011011010100100111101101001011010011000110011110011000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111110011100001110111000100001010000010011100100111101110000011110010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111110100000000100001010010010011011100100001000110010010111101100010001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111110100001000000000101100111001010101011011010000010101000110000010011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111000101111111110110001,
	240'b101100011111111110101011000000000000001101110101110001111011010110101001110001100011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010011111111010101110,
	240'b101011101111111111100000000111110000000000000000001111011000101110100100011100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100111111011111000010011110,
	240'b101100001110111011111111101110010100010000101110001010110010111000110100001011100010111100110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000101111111100010111111111101010110110111,
	240'b110101101100010011111100111111111111100011101101111011011110110111101100111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101111111111111111111011011100000111110111,
	240'b111011101101101111000001111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100000101111001110110111111110,
	240'b111000001111011011011101101001101010001110101010101010111010101010101010101010101010101010101010101010111010101110101011101010111010101010101010101010101010101010101010101010101010101110101011101010011010000110101101111001101111010011110001,
	240'b111010011111110111001001011110001001001110101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101010001000010010001101111010011111110111111010,
	240'b111100001111000010111010110011011110001111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010111101110111000110110010101111110011111111,
	240'b111001001100000011101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100101111111111,
	240'b101110101110001011111111111001101000101101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111001101001011010100110101001101110011100011010011011111010111111111100101111001111,
	240'b101011101111110111110001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001010111110011010100000000000000000000001110001001111111111110101010011110,
	240'b101100001111111110111000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111100101010111000111010000110000110110000000000101000111100001111101110101010,
	240'b101100001111111110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111111111110100110101100001110101100011110000111000011001111000101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111000111101101000110001001001100000010101101100010110111000101111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110110010011001111100010111000010011000111000111001000100110111000011111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101101001001101000000000000000000000000000101111100111011110111111111111110110001,
	240'b101100001111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011011110010101000000010100000010110110110100111010110111111111111110110001,
	240'b101100011111111110100010000000000000000001000000100011011001110010000011011110110110100101000101000111100000000100000000000000000000000000000000000000000000000000000000000011000101011101111000011111100101010100011100111000101111111110110001,
	240'b101100011111111110100000000001111000011011110100111111111111101110000011011010110111101110001101100110001000010101001100000011110000000000000000000000000000000000000000000000000000000000000111000011010000000000011011111000101111111110110001,
	240'b101100011111111110011110011101101111111111111111111111111111111110111101010100010101000101010001010101100110101010001110100101100100111100000110000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111000010111001011111111111111111111111111111111111110111011111000101000001010101010101010101001101010001011000101001000110001001001001010000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111110000111111011111111111111111111111111111111111111111110010010101011001010100010101010101010101010101010100110101001001110100100111010100001000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111111111111111111111111111111111111111111111111111111111111111110111000011001010000010101010101010101010101010101010101010101010001011000011001101001001111000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111111111111111111111111111111111111111111111111111111111111111111101001101011010010101000101010101010101010101010101010101010101010100110101101010011001010011110000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111111111111111111111111111111111111111111111111111111111111111111111110110010001010011110101010101010101010101010101010101010101010101010101001101011011100111010011100000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111111111010111111101111111111111111111111111111111111111111111111111111111111011100010111100101001101010101010101010101010101010101010101010101010101010010011001001001010100010111000000000000000000011100111000101111111110110001,
	240'b101100001111111111100110111110011111111111111111111111111111111111111111111111111111111111111111100110110101000001010101010101010101010101010101010101010101010101010101010100010111101001111001000000100000000000011100111000101111111110110001,
	240'b101100001111111111010001111101001111111111111111111111111111111111111111111111111111111111111111111001010110010001010010010101010101010101010101010101010101010101010101010101010101001110010100001110100000000000011100111000101111111110110001,
	240'b101100011111111110110111110110011111111111111111111111111111111111111111111111111111111111111111111111111010011001010000010101010101010101010101010101010101010101010101010101010101001101100111100010010000010000011011111000101111111110110001,
	240'b101100011111111110100001101010101111111111111111111111111111111111111111111111111111111111111111111111111110110101101011010100100101010101010101010101010101010101010101010101010101010101010010100011110011011000010110111000101111111110110001,
	240'b101100011111111110011011011000111111111011111110111111101111111011111110111111101111111011111110111111101111111110110010010110000101101101011011010110110101101101011011010110110101101101011001011100100111100100011010111000101111111110110001,
	240'b101100011111111110011110001001111001001101000001010000100100001001000010010000100100001001000010010000100100001101000000001010000001110100011101000111010001110100011101000111010001110100011101000111110111001100110111110111111111111110110001,
	240'b101100011111111110100010000000110110111000010010000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000100010001100100110111001111111110110001,
	240'b101100011111111110100010000000000011111001011101000000000000000000000000000000000000000000000000000000000000000000000000000010010000110100000000000000000000000000000000000000000000000000000000000000000001110010000100110111111111111110110001,
	240'b101100001111111110100010000000000000011001110111000111100000000000000000000000000000000000000000000000000000000000000000000000000001000100000011000000000000000000000000000000000000000000000000000000000000010110001110111011001111111010110001,
	240'b101100001111111110100010000000000000000000110010011011110000001000000000000000000000000000000000000000000000000000000000000000000000011100001110000000000000000000000000000000000000000000000000000000000000000010000001111101101111110110110001,
	240'b101100001111111110100010000000000000000000000000011001000100100000000000000000000000000000000000000000000000000000000000000000000000000000010000000001010000000000000000000000000000000000000000000000000000000001101000111110101111110110110001,
	240'b101100001111111110100010000000000000000000000000000011000111101000101011000000000000000000000000000000000000000000000000000000000000000000000110000100000000000000000000000000000000000000000000000000000000000001010011111110011111110110110001,
	240'b101100001111111110100010000000000000000000000000000000000001110101111111001000010000000000000000000000000000000000000000000000000000000000000000000011110000011000000000000000000000000000000000000000000000000001001001111110101111110110110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000100111100000010010100000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000001000111111110101111110110110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000001001001000001000111111000000000000000000000000000000000000000000000000000000000000111000000111000000000000000000000000000000000000000001100001111110111111110110110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000001001101110001011010000001010000000000000000000000000000000000000000000000001100010001000000010000000000000000000000000000010010001110111100001111111010110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000000000000000010010001011000000001010101000101100000000000000000000000000000000000001100000010010000000000000000000000000100111001110100110111101111111110110001,
	240'b101100011111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010010011111100110101100111101000111000000100000000100000100000000000000001110010101110110111000100011111000011111111110110001,
	240'b101100001111111110100001000000110101001101110010010011100001000100000000000000000000000000000000000000000000000000000000000010100011001101011110011101100111101001110101011101110111001101111100010101110000011100011001111000101111111110110001,
	240'b101100001111111110011100001111011111100011000000100001111001010000110010000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100011111001001000010001100001110000000000000000000011100111000101111111110110001,
	240'b101100001111111110011010010101111111111111101010011001110110010110011001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111110011100001110111111000011110111101001100100101101101101011110010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100001111111110100000000100101000110100111000001010100001000100010000011100010001110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111000101111111110110001,
	240'b101100011111111110100001000000000100111101010010000000000000000000000000010100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111000101111111110110001,
	240'b101100011111111110101011000000000000011001101001011001100001111100001011011000110011010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010011111111010101110,
	240'b101011101111111111100000000111110000000000000000001111100111000001111000011000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100111111011111000010011110,
	240'b101100001110111011111111101110010100010000101110001010110011000100111001001100000010111100110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000101111111100010111111111101010110110111,
	240'b110101101100010011111100111111111111100011101101111011011110110111101100111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011011110110111101101111011101111111111111111111011011100000111110111,
	240'b111011101101101111000001111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100000101111001110110111111110,
	240'b111000001111011011011101101001101010001110101010101010111010101010101010101010101010101010101010101010111010101110101011101010111010101010101010101010101010101010101010101010101010101110101011101010011010000110101101111001101111010011110001,
};
assign data = picture[addr];
endmodule