module seaside(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 600;
localparam Y_WIDTH = 430;
parameter [0:1289][2399:0] picture = {
	2400'b110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110010111010100001110110011101110111011101100101010101010101011001100111100010101100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011110111011101110111011101111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111110111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110111011101111111011111110111111101110111111111111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101101111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001011101010000111011101110111011101110110010101010101010101100111100010011011110111101101110111011101110111011101111011101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101111011101110111011101101111011101110111011101110111011101110111011101110111011101110111011101110111011011101111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111110111111111110111011111111111011101110111111101110111111111111111011111111111011101111111011101110111011111111111111101111111111101111111111101111111111111111111111111110111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110010111011101110111010101010011000100001110111011101100110010101000101010101100110100010011011110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001100110111011101110111101110111011101110111011101110111011101110111011101110111011101110111111101111111011101110111011101110111011101110111011101110111011101110110111011110111011101110111011101110111011101110111011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101111111111111111111111111111111111101111111111111110111011111111111011101110111011111111111111111111111111111111111011111110111111101110111011111110111011101110111011101110111111111110111011101110111011101110111011101110111011111111111011101111111011101110111111101111111111101110111111111110111011101111111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110111011011101110111101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110010111010100110011001100110011001100010001000011101100110011001010100010101010110011110011011110111011101110111101101110111101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111101110111011101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111110111111111111111111111111111111111111111111111110111011101110111111111111111011101111111011101111111111101110111011101110111111101110111011101110111011101111111011101110111111111110111111101110111011101110111011101111111111101110111011111110111011111110111111111111111111111111111111101111111011111111111111111110111111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101101110111011101111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b100010101100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001010100110011000100010001000100010001000100001110110011001010100010101010110011110011011110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001100110011001100110011001100110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111111110111111111111111111111111111111111111111111101111111111101110111111101110111011101111111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101111111011111111111111111111111111111111111111101111111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011011110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b010101010110100010101101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110010111011101010101010100110000111011101110111011101110110010101010101010001010110011110001100111011011101110111011101110111011101110111101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110011001100110011001100110011001101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111011111110111011101111111111111111111111111111111111111111111011101111111111111110111011101110111111111111111011111111111111101110111011101110111011101110111011111110111011101110111111101110111011101110111011101110111011111110111011101110111011101110111011101110111011111110111111101110111111111111111111101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b010101010101010101010111101111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001011101111001100101110101001011101110111011001100110011001010101010001010101011010001100110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111111111111111111110111111111111111011101111111011101110111011111110111011111110111111111110111011101111111011101110111011101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b010101010101010001000100010110011100110111011101110111011101110111011101110111011101110111011101110111011101110111001011101110111011110011001011101010000111011001100110010101010101010101000101011010001100110111001101110111011101110111011101110111101101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111111111110111011101110111011101110111011101110111011101111111011101110111011111111111011101110111111101110111011101110111011101110111011101110111011101110111011101110111111101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b010101010100010001010101010001010111101111011101110111011101110111011101110111011101110111011101110111011101110111011100101110111010101010101010101110101001011101100101010101010101010101010100011010001011101110101101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110110111011110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011111110111011101110111011111111111011101110111011101111111111101110111011101110111011101110111011101111111011101110111011101110111011101111111111101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b010101010101010001000100010001000101011010101101110111011101110111001101110111011101110111011101110111011101110111011101110111001011101010011010101010101001100101110110010101010100010101010100010101111010100110101100110111011101110111011110111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111110111011101110111011101110111111101110111111111110111011101110111011101111111111111110111011111111111111111111111111111111111111111110111011101110111011111110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b010101010101010101010101010001000100010001011001110111011101110110111100110011011101110111011101110111011101110111011101110111011101110010111001100010011001100110000111010101010100010001010100010101111000100010101011110111011101110111011110111011011110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111111101110111111101110111011101110111011101110111011101110111111101110111011101111111011111111111111111111111111101111111011101110111011101110111011101110111011101111111111111110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b011001100101010101010101010101000100010001000101100011001101110110111011101111001101110111011101110111011101110111011101110111011101110111001010100110001000100010000111011001010100010001000100010101100111100010101100110111011101110111011101110111101110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011111110111011101110111011101110111111111111111011101111111111101111111011111110111011101110111111101111111111111110111011111111111111111111111111111110111111111110111011101110111011101110111011101111111011101110111011101111111011101111111011101110111011101110111011101110111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b011101100110011001100101010101010101010101010101010101111010110010111001101010101100110111011101110111011101110111011101110111011101110111001010100110000111011101110111011001100100010001000100010101100111100010101100110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111001101110011001100110011001100110011001100110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111110111111111111111011101110111011101110111011101110111011101110111011111110111011111111111011111110111111111110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b100110000111011101100110010101010101010101010101010101010110100010101000100010101011110111011101110111011101110111011101110111011100110010111011101010011000011101110110011001010101010001000100010001100111100010101011110111011101110111011101110111011101111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011101110111011101110111011101110111011101110111011011110111011101110111011101110111011101110111111101110111011101111111111101110111011101110111111111111111111111110111111101110111011111110111011101110111011101110111111101110111011101111111011111111111111111111111011111111111011101110111011101110111011111110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101010011001100001110110011001100101010101010101010101010101010101110111011110011001101111001101110111011101110111011101110111001011101110111011101010011000011101100110011001010101010101000100010001010111100110101010110011011101110111011101110111101110110111101110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011100110011001100110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011110111011101101111011011110111011101110111011101110111011101110111011101110111011101111111011101110111111111110111011101111111011101110111111101110111011101110111111101110111011101110111011101110111011101111111011101111111011111111111111111111111111101110111111101110111011101110111011101110111111101110111011101111111111101111111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101010101001100001110111011001100110010101010101010101010101010101010110011101111000100110111100110111011101110111011100110011001011101110011001101010101001100001110110010101010100010101000100010001010111100110011010110011011101110111011101110111011110111011101110110111101101111011101110111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110111011101110111011101110111111101110111011101110111011101110111011101111111111111110111011101111111011101111111011111111111011101110111011101111111011101110111011101110111011101110111111101110111011101110111111101111111111111111111111111111111111111111111011111110111011101110111011101111111011101110111011111111111011101111111111101110111011101110111011101110111011101111111111101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101010101001100001110111011101100110011001100101010101010101010101010101010101100111100010011010110011011101110111011100110010111010100110011001100010011001100101110110010101010100010001000100010001010110011110001010101111011101110111011101110111101110110111101110110111011110110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011110111011101101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101110111011101110111111101110111111101110111011101110111011101110111111111110111011101110111011101110111011111110111011101110111011101110111011101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111101110111011111111111011111110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101010011000100010001000100010011001100001110110010101010101010001000101010101010110100010001001101011001101110111011100110010111010100110001000100010001000100010010111010101000100010001010100010001000110011010001001101010111100110111011101110111011101111011011101111011101110110111011110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011110111011101110111011101110111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101110111111101110111011101110111011111110111111111110111011101111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111101110111111111111111111111111111111111111111111101111111111101110111011101110111011101110111111101111111011101111111111101110111011111111111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b100101111000100010001001101010101011101010011000011101100101010101010100010001010101011110001000100110101100110011011101110010111010100110001000011101110111011110001000011001010100010001000101010001000101011010001000101010101011110111011101110111011101111011011101110111101110111011011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101111111111101110111011111111111011101111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111110111111111111111111111111111111101110111011101110111011101111111111101111111111101111111011101110111111111110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b100010001001100010001000100010001000011101111000100001110110010101000100010001000101011001111000100010001010101111001101110111001011100110000111011101110110011001110111011101100100010001000101010101000101011001111000100110011010110111011101110111011101110111011101110111011101111011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111101110111011101111111011111111111111101111111111111110111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111111110111111111111111011111111111111101111111111111110111011101111111111111111111011101110111011111111111011111111111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b100110000111011110000111011001010101010101000100010101100101010101000100010001000101010101100111011110001000101011001100110011001011101010101000011101100110010101010110011101110101010001000101010101000100010101101000100010001011110111011101110111011101110111011101110111011101110111011101111011101110110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111111101110111011101111111111101110111011111110111011111111111111101110111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111011101111111111111111111011101111111111101110111011111110111111101111111111111111111111101110111011111111111111111110111011111110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110110111011101110111011101110111011101110111011101110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b100110011010101110101001100001110101010001000100010001000101010101010101010101010101010101010110011101110111100010101011110011001100101110101001100101110110010101010101011001100110010101000101010101010100010001100111100010001011110011011101110111011101110111011101110111011101110111011101110111011101110111001100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111111111111111111111111111111111111111011101111111011101111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011111111111111111111111111101110111111111111111011111110111011101110111111111110111111101110111111111111111111111110111011101111111111101110111011111111111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011101101111011011101110111011101110111011101110111011101110111011100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b110011001100101110101010100110011000011101010100010000110011010001000101010101010101010101010101011001100111011110001001101111001011101110101001100010000111011001000100010001010101011001010101010101010100001101010111100010001010101111001101110111011101110111011101110111011101110111011101110111011101110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111011101111111111101110111111101111111011111111111111111110111011101110111011111111111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111110111011101111111111111111111011111110111111111111111111101110111111101110111111111111111011101110111011111111111111101110111111101110111111101110111011101111111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110110111011101110111011101110111011101110111011101110111011100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b110011001011101010011000100010001000100010000111010101000011001101000100010101100110011001010100010101100110011101111000100110011001100110101010100101110111011101100100010001000100010101100110010101000100001101010111011110011001101111001101110011011101110111011101110111011101110111011101110010111011101111001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101111111111101110111011101110111011101110111111111110111111111111111111101110111011111111111111101110111011101111111111101110111111111110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101111111111111111111111111111111011111110111111111110111111111110111111111111111111101110111111111110111111111110111011101111111111111110111011101110111011101110111011101110111111101111111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101110101001100110001000011101111000100010011000011001010011001100110011010001010110011001010101010101010101011001100111011101110111100110011001100110000110011001100101010000110100010001010101010101000011001101010110100010001000101010111100110011011101110111011101110111011101110111011101101010001001100110011010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111111101110111011111111111011101110111011101111111111111111111111111111111111101110111011101111111011101110111011101110111011101110111011101110111011111111111011101110111011101111111111111110111111111111111111101111111111111110111011111110111111111111111111111111111111111110111011101110111111101110111011101110111111101110111011101110111011101110111011101110111011101110111111101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110110111011101110111011101110111011101110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101110111010101010011000011101110111011101111000011101100101001100110011010001010110011001100110010101010101010101100110011001100110011001110111011101110111011001010110010101000011001101000100010101000011001101000111100010001000100010101011110011011101110111011101110111011101110111011011100001100110011001101000101111011101111011101110111011101110111011101110111011101110111011101110111011101101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111110111011111111111111111111111111101110111011101110111111111111111011101110111011101110111011111110111011101110111011101110111011101110111011111110111111111110111011101111111011101111111111111111111011111110111111111111111111101111111111111111111011111110111111111110111011101111111111111111111011101110111011101110111011101110111011111110111011111110111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100101110111100110011001101110111011101110111011101110111011101110111011101110111011101110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101,
	2400'b101110111011101010101010100110011000100010001000011101100101010101000011001100110101011001110110010101010101011001010101010101100110011001100110011001110110011001010101010101010011001100110100010001000011001101000111100001110111100010011011110011001101110111011101110111011101110010111000010101000101010101111010101110111100110111011101111011101110110111011101110111011101110111101101110010111100110011011101110011001100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111101110111111111111111111111111111011101110111011101111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111111111110111011101110111111101111111011101110111011101111111111111110111011101111111111111111111111101110111011101110111111111111111111111110111011101111111011101110111011101110111011101111111011101110111111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111101101111011011101110111011101110111011101110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100101110111100110011001101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111001100,
	2400'b110011001011101010101010100110011000100110001001100010000110010101000011001100100011010001100110010101010101011001100101010101010101010101100110011001100110010101010101010001010101001100110100010000110011001101000111100001110111100010011011101111001100110011011100110011001011101010000101010001000100011001110111011110001000100110101011110111011110110111011101110111011101110111011011101010111101110111001011101010111100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111110111111101110111011101111111011111111111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011111111111111111111111111111111111011101110111011111111111111111111111011101111111111111111111011101110111111101110111111111111111111101110111111101111111011111110111011101111111111101111111011101111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101111011011101110111011101110111011101110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100101111001100110011001100110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001101110111001101110111011101110111011101110111011101110111001101110111001100,
	2400'b110011001100110010111011101010011000100001111000011101100101010101000011001100100010001101010101010101010100010101100110010101010101010001010110011001100101010101010100010101000101010101000011001100110010001101000110011101110111011110011010101111001100110011001100101110101001011101100100010001000101010101100111011101111000100010011001101010111100110111011101110111101101110010011010110011011100101010101011110011001100110011001100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111111101111111111111111111111111110111011101111111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111011101111111111111111111111101110111011111110111011101111111111111111111011111111111111101111111111111110111011101111111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111101110111011101110110111011101110111001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100101110111100110011001100110011001101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111001100110011001100110111001100,
	2400'b110011001011101110111011101010101010100001110101010101010101010001000011001100100010001001000101010101010100010001010110011001010100010101010101010101100110010101010100010001000100010001010011001100110010001101010110011101100111100010001001101110111100101110111010100101110110010101000100010001010110011001100110011101111000100010001001100110011001101010111100110011001010100010101101110010101010101010111010100110011000100001110111011101111000100010011010101111001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111111111111111111101110111011111111111011101111111011111110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111111111111111111101111111111101110111011101110111011101110111111111111111011111111111111101111111111111110111011101111111011101111111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101111011101101111011101110111011011101110111011101110111011101110111001100110111011100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110010111011101111001100110011001100110111011101110111001100110011001011101111001100101111001100110011001100110011001100110011011101110111011101110111011101110111011100110011001100110011001100,
	2400'b110011001100110010111010101010101001100001100101010001000100010001000100001100100010001000110101010101010101010001000101010101010101010101000100010001100110011001010100010000110011010001000100001100110010001101000110011101100110100001111000100110111011100110010111011001010101010001000100011001110111011001100111011101111000100010001000100110011001101010101010101001110110100010111000011001010110011001100110011001100101010101100110011001100110011101111000100010001001101111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101111111011101110111111111110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111011101111111111111110111011111110111111111110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111011101110111011101111111011101111111111101110111111111111111011111111111111101111111111101111111111101110111011101110111011111111111011111110111111101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001011101110111011101110111011110011001100110011011101110111001100110010111011101110111011101110111011110011001100110011001100110011001100110011001100110011011101110111011100110011001100110011001100,
	2400'b110111001100110011001011101110101010100110000111010101000011001100110100010001000011001000100100010101010101010001000100010101000101010101010101010001000110011001010100010000110011010001000100010000100010001101000101011001100110010101010111100110101001100001110101010001000100010001010110011101100110011001100111011101111000100010001001100010001000100110000110010101000100010101010100010001010100010101100110011101100110011001100110011001100110011001110111100010001000100110101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111011101111111111111111111011111110111111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111110111011101111111011101111111111101110111111111111111011101111111011111111111111111111111111101110111111101110111111111110111011111110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001011101110111011101110111011110011001100110011011101110011001100110010111011101110111011101110111011101110111011110011001100110011001100110011001100110011011101110011001100110011001100110010111011,
	2400'b110111011101110111011100110010111010100110011000011101100100001100110011001100110011001100100011010101010101010001000100010001010100010001000100010101010101010101010100010000110011001100110100010000110010001101000101011001010110010001010110100010000111011001010100010001000100010101100101011001100111100010001000100110011001100110011001100110000111011001000011001100110011001101000100010101100111011001100110011110001000011101110111011101110111011101110111011101111000100110011011110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011111111111111101111111111111111111011111111111111111110111111101111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011111110111011101110111111111111111111111111111111111111111111101110111111101110111111101110111111101111111011111111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011011100110011001100101110111011101110111011101110111011110011001100110011011100110011001100101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001011101110111011,
	2400'b110111011101110011001100110010111010100110001000100001110110010101000011001000100010001100110011010001010101010101000100010001010101010001000011010001010101010001000100010000110011001100110100010000110010001101000101010101010100010001000101011001110110010001000100001101000101010101010101011001111000100010011001100110011001100110011000100001100100001100110011001100110011010001000101011001111000100010000111011001100111100010000111100110101010101010011000011101110111011110001001101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011111111111111101111111111111110111011111111111011111111111111101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111101110111011111110111011111111111111111111111111111111111011101110111011111111111111111110111111101111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001011101110111011101110111011101110111011101111001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100101110111011101110111011,
	2400'b100110111100110011001011101110111010101010011001100001110111011001010100001100100010001000100010001101000101010101000100010001000011001100110100001101000100010000110011010000110011001100110011001100110010001101000100010101000011010001000100010101100101010001000100010001000100010001010110011101111000100010001000100010011001100110000110010100110011001000110011001100110100010001010110011001111000100010001000011101100110011110001000100010101011110011001011100110000111011101110111100010011100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101111111111111110111111111111111011101110111011101111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111011101110111011101110111011111111111011101110111111101110111111111110111111101110111011101111111111111110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001011101110111011101110111011101110111011101110111100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001011101110111011101110111011,
	2400'b010001101010110011001011101110101010101010101001100010000111011101100101010000100010001000100010001000110100010101010101010001000100001100110011001100110011001100110010001100110011001100110011001100110010001101000100010000110011001101000100010001000100010001000100010001000101010101100110011101110111100010011000100010001000011101010011001000100010001100110011001100110100010001010101011001111000100010001000100001110110011110001000100010001011110111101101110010101001100001110111011101111000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111110111011101111111011101110111011101110111011111110111011101110111011101110111011101110111111101111111011111111111111111111111111111110111011101110111011101111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101111111011111111111111101110111111101110111111111110111111101110111111111111111111111110111011101110111011101111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111001101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110010111011101110111011101110111011,
	2400'b001100110101100010111100101110101001100110101001100110001000011101100110010101000011001000100001000100100011010001010101010001000101010000110011001101000011001100110010001000100011001100100010001000100010001100110100010000110011001100110100010001000100010001000100010001010101010101100111011110001001100110011001100001110101001100110010001000110011001100110100010001010101010101010101010101100111100010011001100010000111011101111000100110001001101111011101110111011011101010001000011101110111100111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111110111011101110111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011111111111111111110111111111110111011111111111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011111111111111101110111011101111111111101110111011111110111111111111111111111111111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110110111011101110111011101110111011101110111011101110111001100110011001100110011011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001011101110111011101110111011101110111011,
	2400'b001000100010010001111001101010101010101010011001100110011000100001110110010101000100001100100010000100010010001101000100010001000101010000110011001100110011001100110010001000100010001000100010001000100010001100110100001100110011001100110011010001000011001101000100010101000101010101100110011110001001100110011000011101010011001000100011001100110011001100110100010101100110011001010101010101100110011110001001100110011000011101111000100110011000100111001101111011101101110110101000100001110110011110101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111110111011101110111111101110111011101110111011111110111011101110111011101110111011101110111011101111111011101110111111111110111011101110111111101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101111111011101111111011101111111111111110111011101111111111101111111011101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011100110011001100110011001100110011001101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101110111011101110111011101110111011101110111011,
	2400'b001100100010001000110101011110011010101010101001100110011000011101110111011101010100001100100001000100010001001000110011010001000100010101010011001100100010001100110010001000100010001000100010001000100010001100110100001100110011001100110011001100110011001100110100010001000101010101100111011110001000100010000111010000110010001000110011001101000100010001000100010001010111011101100110011001100110011101111000100110101001100010001000100110111001100110101101111011101110111011001010100101110111011101111010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011111111111111101110111111101111111111111110111011101110111111101110111011111110111111101110111111111111111111111111111111111110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101111111011111111111011111110111011101111111111111111111011101110111111111111111011101110111011111110111011111110111011111110111011101111111011101110111011101110111011111110111011101110111111101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110111011101110011001100110011001100110011001100110011001100110011001011110011001100110011001011101110111011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100101110111011101110111011101110111011101110111011,
	2400'b001100100010001000100010001101010111100110011001100110001000011101110110011001000100001100100010000100010001001000100011010001000100010101010100001100100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001101000100010001010101010101100111011101111000011101100100001100100011001101000100010001000100010101010101010001000101011101110111011101110111011101111000100110101010100110001000100110111100101010011011110111101110111011101101101110000111011101111000101111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101111111111101110111011111111111111101110111011101111111111101110111011101110111011101110111011111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011111111111011111111111111111111111111111111111011101110111011111111111011101111111111101111111011111110111011111110111011101110111011101110111011111110111111101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011011100110011001100110011001100110011001100110011001100101111001100110011001100110011001100101111001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100101110111011101110111011101110111011101110111011,
	2400'b010000110010001000100010001000100011010101111001100110001000100001110110010101010100010000110010000100010001000100100010001101000100010001010101010000100010001000010010001000100010001000100010001000100010001000110011001100110011001100110011001100110011010000110100010101010101010101010101011001110111011001000010001100110100010001000100010001010101010101010101010101010101011001111000100010001000100010001000100110101010101010011000100010101100110010101010110011101110111011101110110110111000100010000111100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111111111110111011101110111011111110111011101110111011101110111011101110111011101110111111101110111011101110111111111111111111111111111011101111111111101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111011111111111011111110111111111111111111111110111011101111111111111111111011111111111111101111111111111110111011111110111011101110111011101111111111111111111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011110011001100110011001100110011001100110011001100101111001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110010111011101110111011101110111011101110111011,
	2400'b010001000011001000100010001000100010001101000101011010001000011101100110011001100101010000110010001000010001000100010001001000110011010001010101010100110010000100010001001000100010001000100010001000100010001000110100001100110011001100110011001100110011001101000100010001000100010001010101010101100101010000100010001100110011010001000100010101010101010101010110011001010110011001111000100010011001100110011001100110011010101010101010100110011011110111011011101011011110111011101110111011101011101110101000011110011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111111111110111111101110111111101110111011101110111011101110111011101110111011101110111011111110111011101110111111101111111111111111111111111110111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101111111111111111111111111110111011101111111111111111111011111111111011111111111111101110111111101110111011101110111011101110111111101111111111101111111111101111111011101110111011101110111111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100101110111011110011001100110010111100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110010111011101110111011110011001100110011001011,
	2400'b010001000011001100100010001000100010001000110010001101000100011001100110011001010101010101010100001100100001000100010001001000100011001101000101010101000010000100010001000100010010001000100010001000100010001100110011001101000011001100110011001100110100001100110011001100110100010001000100010101010100001100100011001100110011010001000101010101100110011001100110011101100110011001111000100010011011101010101010101010101010101110111011101010011010110011011101101111001110111011101110111011101110110111011011100010001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101110111111101110111011111110111111111110111011101110111111101111111011101110111011101110111011101110111011101111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101111111111111111111111111110111011101111111111101111111111111111111111111111111111111111111111111111111011101110111011111111111111101111111111101111111111111111111011101110111011101110111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110010111011101111001100110011001100110011001100,
	2400'b001000100010001000100010001000100010001000010010001000100010001000110101010101010110011001110111010100110010000100010001000100010010001100110100010101010011001000010001000100010001001000100010001000100010010001000011010000110011001100110011001100110011001100110011001101000100010001000101010100110010001100110011010001000100010001000101010101100110011101100110011101110110011001111000100110011010110010111011101110111010101011001100101110111010101111001101110111001101111011101110111011101110111011101101101110011001110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011111110111011101111111011101110111011101110111111101110111011111111111011101111111111111111111111111111111111111111111111111110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111101111111011111111111111111111111111111111111111101111111111101110111011101111111011101110111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100,
	2400'b001000100010000100100010001000100010001000010010001000100010000100010011011001100110011101100101010000110011001000010001000100010001001000100011001101000011001000010001000100010001000100100010001000100011001100110011001100110011001100110011001100100011001100110011001100110100010001000100001100100010001100110011010001000100010001000100010101100110100010000111011101110111011001101000100110011010101111011100110011001011101111001101110011001011101111001101110111011101111011101110111011101110111011101110111011001010101011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111101110111011111110111011101110111111101110111011101111111111101110111011101110111011101111111111101111111111111111111111101111111111101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111110111111111110111011111111111111111111111011111111111111111111111111111110111111101110111011101111111111111111111111111111111111101110111011101110111011101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110010111100101110111011110011001100110011001100110011001100110010111100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100101111001100110011001100110011001100,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001101000110011101100101010101000010001000010001000100010001000100010010001000100010001000010001000100010001000100100010001000100010001100110010001100110010001000110010001100110011001100110011001100110011001100110011001000100011001100110011001100110100010001000100010101100111011110000111011101110111011101110111100110011001101011001101110111011100110010111101110111011101101111001101110111011101110111101110111011101110111011101110111011101101101111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101110111111111110111011101110111011101110111011101110111011101111111011111111111011101110111011101110111011101111111111101111111111111111111111101111111111111111111111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111011111111111111101111111111111111111011111111111111111111111111111111111111111110111011101110111111111111111011101111111111111111111111111110111011101111111111101110111011111111111111101111111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001100110011001100110111011101110111011101111011101110111011101110111011101110111011101110111011101110110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111001100110011001100101111001100110011001100110011001100110011001100110011001100110010111011101110111100110011001100110011001100110011001100110010111100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100,
	2400'b001000100010001000100010001000100010001000110010001000100010001000110010000100010011011001100101010001000011001000010001000100010001000100010001000100010001001000100010000100010001000100100010001000100010001000100010001000100011001000100011001100100010001000100010001100110011001100100010001000110011001101000011001100110100010001000100010101100111100010001000011101110111100010001000100110011010101010111100110111011101110111001101111011101110110111001101111011101110111011101110111011101110111011101110111011101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111011111111111011111111111011111110111011101110111111101110111011101110111111111111111111111111111111101111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111110111011111111111111101110111011111111111111111111111111111110111111111110111111111111111111111111111011101111111111101111111111111110111011101110111011101110111111111110111011111110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110011001101110111101110111011101110111011101110111011101110111011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101101111011101101110111011101110111011101110111011101110111001011101110111011101110111011110011001100101111001100110011001100110011001011101111001100101110111100110011001100110011001100110011001100110011001011101110111100101110111100110010111011101110111011101110111011101110111011101110111011101110111011101010011001011101111000100110101010101110111100110011001100110011001100110011001100101110111011110011001100110011001100,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010000100010001001001000100010000110010001000100001000100010001000100010001000100010001000100100010001000010010000100100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000100010001000100010001010111100010001000100010001000100010011010100110111010101010111011110111101101110111011101111011101110111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111101110111011101110111011101110111011111110111111101110111111101110111011101111111111111111111111111111111011111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111011111110111111111111111011101111111111111110111111111111111011101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110011001100110011001100110011001100110111101110111011101110111011101110111011101110110111011101110011001100110011011101111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110011001100101110111011101110111011101110111011101110111100101111001100110011001011101110111011101110111100110011001100110011001100110011001100110010111100101110111011101110111100110010111011101110111011101110111011101110111011101110111011101110111011100101110110011001111000101010101011101110111100110011001100110011001100110011001100101110111011110011001100110011001100,
	2400'b001000100010001000100010000100010010001000100010001000100010001000100010001000010001000100010010001000100010001000100010000100010001000100010001000100010001000100010010001000100010000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011010000110011001100110011010001000100010101010110011101111000100110011001100110011010101010101011101010111100110011011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111111110111111101110111111111111111111111111111111111110111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111111111111011101110111011101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111101110111111111110111111101111111011111110111111111110111111111110111011101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011011101110111001100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110011001100110011001100110011001100110011011110111011101110111011101110111011011101110011001100110011001100110011011101111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011100110010111011101110111011101110111011101110111011110010111011110010111011101110111011101110111011101110111011101110111100110011001100110011001100101110111011101110111011101110111100110010111011101110111011101110111011101110111011101110111011101110111001011001010101100010011010101010111011101110111100110011001100110011001100110011001100101110111011110011001100110011001100,
	2400'b001000100010001000100010000100010001000100010001000100010001000100010010001000010001000100010001000100100001000100010001000100010001000100010001000100010001000100010001000100100010001000010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000110011001100110100001101000100010001000101010101010110011101111000100110101010101010101010101111001100110010111100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111101110111011101111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101111111011111110111011101110111011111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111110111011101111111111111111111111111111111111101110111011111110111111111110111011111110111011101111111011101110111011101111111111101110111011101110111011101110111011101111111111101101110111001100110011001100110011001100110111101110111011101110111011011101110111101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110010111100110011001100110011001100110011011101111011101110111011101110111011011100110011001100110011001100110011001101110111011101110111011110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011110011001011110010111011101110111011110010111011110011001100110011001011101110111011101110111011101110111011101110111011101010010101010001100111011110001000100110101011101111001100110011001100110011001100110011001100101110111011110011001100110011001100,
	2400'b001100110010001000100010001000010001001000010001000100010001001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100100011001100110100010001000100010001000101010101100110011110001000100010101011101010101011101111011101110011001100110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101111111111101111111011101110111111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111111101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111111111111111111111111111011101111111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111101110111111111111111111101110111111111110111011101111111011111111111111111111111011101110111111101110111011101110111011101111111111101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110111101110111011101101110111001100110111011101110111011110111011101110111011101110111011101110111011101101110111001100110011001100110011001011101110111100110011001100110011001101111011101110111011101110110111001100110011001100110011001100110011001100110011001100110011001101110111101110111011101110111011101101110111011101110111011101110111001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011101111001011101111001100110010111011101111001100101111001100110011001100110011001011101110111011101110111011101110111011101110101001100101010100010101100111011110001000100110011010101111001100110011001100110011001100110011001100110011001100110011001100110011001100,
	2400'b010001000011001100110010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100011001100110011001100110011001100100010001100110011001100110100010001000100010101010101011001100111011110001001100110011010101110101010110011011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101111111111111111111011111111111111111110111111111111111111101111111111111111111111111111111111111111111111111111111011101111111011101110111011101110111011101110111011111110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111111111111111011111110111111111111111111111111111111111111111011111110111011111111111111111111111111111111111111111111111111111111111011101110111111111111111111101110111111111110111011111110111011111111111111111110111011111110111111101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110011001100110011001101111011101110111011011100110011001100110011001100110111011101111011101110111011101110111011101110111011011101110011001100110011001100101110111011101110111011110011001100110011001101111011101110111011101101110111001100110011001100110011001100110011001100110011001100110011001100110111011110111011101110111011011101110111011101110111011101110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111100101111001100101111001100110010111011101111001100110011001100110011001100110011001011101110111011101110111011101110111011100101100110011001000101011001100111011110001000100010011010101111001100110011001100110011001100110011001100110011001100110011001100101110111011,
	2400'b010101010100010000110010001000100010001000010001000100100001001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010000100010001000100100010001000100010001000100010001000100010001100110011001100110100010001000100001100100010001000110011001100110100010001000100010001010101011001110111100001111000101010101010101111001010101111011110111011011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011111110111111101111111111101111111011111111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101111111111101111111111111110111011101111111111111111111111111111111111111110111111111111111111111111111111111110111111111111111111111111111111111111111011111111111111111111111011111111111111111110111011111111111011111111111111111110111011101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110110111001100110011001100110011001100110011011110111011101110110111001100110011001100110011001100110011011101111011101110111011101110111011101110111011011100110011001100110011001011101110111011101110111011110011001100110011001101110111101110111011101101110011001100110011001100110011001100110011001100110011001100110011001100110011011110111011101110111011011101110111011101110111011100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011101110111011110011001100110011001011101111001100110011001100110011001100110011001100110011001011101110111011101110111011101110111001011001000100010001000110011001100110011101111000100110101011101111001100110011001100110011001100110011001100110011001100110011001100101110111011,
	2400'b011001100110010101000100010001000011001000010001001000100001001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100001000100010001001000100010001000100010001000100010001000100010001100110011001100110011001000100010001000110011001100110100010001000100010001000101010101100111100010001000100110111010101111001100101111001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111101111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101111111011101111111111101111111111111110111111111111111111101111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111110111111111111111011111111111111111111111011101111111111101110111011101110111011101101110111101110111011101110111011101110111011101110110111001100110011001100110011001100110011011110111011101101110011001100110011001100110011001100110011001101111011101110111011101110111011011110110111011100110011001100110010111011101110111011101110111011101111001100110011001100110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011011110111011101110110111011101110111011101110111001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001011101110111100110011001100110011001100110011001100110011001011101110111011101110111011101110010101001100110011001101000111011001100111011101111000100110101011110011001100110011001100110011001100110011001100110011001100110011001100101110111011,
	2400'b011101111000011101100110011001010011001000100010001000100001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001100110011010001000100010101000101010001000101010101010110100110101001100010011100101111001101110111001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101111111111111110111011101110111011101111111111111111111111111111111111111111111111111111111111101110111111101110111011101111111111111110111111111111111111111111111011101110111011111111111011101110111011101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101111111111111111111111111110111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111011101111111011101110111011111111111011011101110111101110110111011101110111011110111011101110111011101110111011101101110111001100110011001100110011001100110111011101110111001100110011001100110011001100110011001100110011001101111011101110111011101101110111011110110111011100110011001100101110111011101110111011101110111011101110111100110011001100110011001101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101111011101110110111011101110111011101110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100101110111100110011001100110011001100110011001100110011001100110011001011101110111011101110111011100101010100001100110011001101010111011001100110011110001000100110101011101111001100110011001100110011001100110011001100110011001100110011001100110010111011,
	2400'b100010011000100010001000100001010011010000110010001000100001001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001000100010101010110011001010101010101010101100010111011101010011010110111001101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101110111011101110111011101111111011111110111011111110111011101111111111111111111111101111111111111111111111111111111111101110111011101110111011101110111111111110111111111111111111101111111111101111111011101110111011101110111011101110111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111101111111111111110111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111110111011101110111111111110110111011100110111011101110011001100110111011110111011101110111011101110111011101101110111001100110011001100110011001100110011011101110011001100110011001100110011001100110011001100110011001101110111011101110111011100110011011101110011001100110011001011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110010111100110011001100110011001100110011001100110011001100110010111011101110111011101110111010011001000011001100110011010001100111011001100110011101111000100110101011101111001100110011001100110011001100110011001100110011001100110011001100110010111011,
	2400'b100110011001101010101001011101000101010101000100001100100010001000100001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001000100010101110110011101110111011001100101011110101100110010111010110011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111111111110111111111110111111111111111111111111111011111111111111111111111111111111111111101110111111111111111011101110111111101110111111101111111111101111111111111111111011101110111011101111111111101110111011101111111111101110111111101110111011101110111011101110111011101110111011101111111011101110111011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111011101110111111101111111111101101110111001100110011001100110011001100110111011110111011101110111011101110111011011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110010111011101110111100101111001100110011001100110011001100101110111011101110111011101110111001010101000011001100110011010101110111011001100110011110001000100110101011110011001100110011001100110011001100110011001100110011001100110011001100110010111011,
	2400'b100110011010101010101001011001010111010101000110010100110010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001001000100001001000100010000100100010001000100010001000100010001000100010001000100011001100110011001000100010001000100010001000110011001100110100010001010101010101100111011001111000100101110110011110011011110111001100110011011110110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101111111111101110111011101110111011101111111111111110111011101110111111111111111111111111111111111111111111111111111111101110111111101110111011111111111011111110111111111110111011101110111111101111111111101111111011101110111011111111111011101110111111101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111101110111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011111111111011011101110011001100110011001100110011001100110111011110111011101110111011101110110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011100110011001100110011001100101110111100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110010111100101110111011101111001100110011001100110011001011101110111011101110111011101110100111010000110011001100110011010110000111011001100110011101111000100110101011110011001100110011001100110011001100110011001100110011001100110011001100101110111011,
	2400'b100010011010101010011000010101110111010001100111011001000100001100100011001000100010000100010001000100010001000100010001000100010001000100010001000100010001001000100010000100100010001000010010001000100010001000100010001000100010001000100010001100110011001100110010001000100010001100110011001101000100010001000110011001010110011101101000101010010111011110001010110111011100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111111101110111011101110111011101110111011101110111011101110111011101111111111101111111011111111111111111111111111111111111111111111111111111110111011111111111011101110111011111111111011111111111111101110111111111111111011101110111011111111111111101110111011101110111111111110111011101110111111111111111111111110111111101110111011101110111111101110111011101110111011101110111111101110111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111011101110111011101110110111011101110011011100110011001100110011001100110111011110111011101110111011101110110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111001100110011001100110011001100101110111011101111001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110010111011101110111011101111001100110011001100110010111011101110111011101110111011101010100111010000110011001100110011010001110111011001100110011101111000100110111011110011001100110011001100110011001100110011001100110011001100110010111011101110111011,
	2400'b100110011001100110010110011001110110011010000111011001100110010001000011001000010010001000100001000100010001000100010001000100010001000100010001000100010001001000100010000100100010001000100010001000100010001000100010001000100010001000100010001100110011001100110010001000100010001100110011001101000100010101010101011101110101011001110111100110101000100010011001110011011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101111111111101111111111101111111111101111111011111111111111111111111111111110111111111111111011111111111011111110111011101111111111111110111111111111111011101111111011111111111111111110111111111110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111110111111111110111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111011101110111001100110011001100110011001100110111011110111011101110111011101110110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001011110011001100101111001100110010111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110011001100110011001100110011001011101110111011101110111011101111001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111010101010101011101110111011101110111011101110111100110011001100110010111011101110111011101110111010100110010111010100110011001100110011010001100111011001100110011001111000101010111011101111001100110011001100110011001100101111001100101110111011101110111011101110111011,
	2400'b100110011001100101110111011101110110011110000110011101100101010001010100001000010001001000100001000100010001000100100001000100010001000100010001000100010001000100100010001000100001000100100010001000100010001000100010001000100010001000100010001100110010001000100010001000100010001100110011001100110100010001010101010101110111011001110111100010011001011110011010101011001101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101111111111111110111011101110111011111110111011111111111011101110111011111110111111101111111111111110111011111110111011101111111011101111111111101110111111111111111111111111111011111110111011101110111011101111111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111110111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110110111011101110111011100110011001100110011001100110111011101110111101110111011101101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111010100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110000110010000110011001100110011010001100111011001100110011110001001101010101011101111001100110011001100110011001011101110111011101110111011101110111011101110111011,
	2400'b101010011001100110001000100001110111100001110111011001100110010101000011001000100010001000100010000100010001000100010010000100010001000100010001000100010001000100100010001000100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001000100010001000101010101010111011101111001100010001010101111001101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011101110111011111110111111111111111111111111111011111111111111101111111111111110111011101110111011101110111011111111111111111111111111111111111111111110111111111111111011101110111111111110111011101110111011101110111011101111111111101110111011101111111011101110111011111110111011101111111111111110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110111011101110111011101110111001100110011001100110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111010100110001000100110101011101110111011101110111011101110111011101110111011101110111011101010011001100001110110010000110011001100110011010001100111011001100110011110001001101010111011101111001100110011001100110010111011101110111011101010101011101110111011101110111011,
	2400'b100010001001100110011010100110001000100010000111011001100110010101000100001100100011001000100010000100100010001000100010001000010001000100010001000100010001000100010010001100110010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000110010001000100010001100110100001100110100010001000101011001100111100010001010101011001101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011111111111111101110111011111110111011101110111011101111111011111111111011101110111011101111111111111111111111111111111111111111111111101111111011101110111011101110111111111111111111111111111111111111111111101111111111111111111111111111111111101110111111111110111011111111111011101110111011101110111011101110111111111111111011101110111011101111111111111110111011101111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110110111011101110111011101110011001100110011001100110011011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110010111100110011001100101111001100101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010001000100010001010101110111011101110111011101110111011101110111011101110111010101010011000011101100101010000110011001100110011010001010110010101100111011110001000100110111011101110111100110011001100110010111011101110101010101010101010101010111011101110111011,
	2400'b001101000101011001101000100010000111100010000111011101110110011001100110010101010100001000100010001000100010001000100010001000100001000100010001000100010001000100010001001101010100001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100011001100110011001100110100010001010101011001111000100110111100110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101111111111111110111011101110111011101111111011101110111011101110111111111111111111101110111011101111111011101111111011111111111111111110111011101110111011101110111011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110111011101110111011101110111011111111111011101111111111101110111011101110111011111111111111111110111111111111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111111111111111111111111111111111011101101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110010111011110011001011101111001100110011001100110011001100110011001100110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010111011110001000101010111011101110111011101110111011101110111011101110111010100110011000011101100101010000110011001100110011010001010101010101100111011110001000100110101011101110111011101111001011101110111010101010011001101010101010101010101010101110101011,
	2400'b000100010010001000100011010000110011001101000101011001100111100010000111011101100100001100110010001000110011001000100010001000100010000100010001000100010001001000100001001001000110010100110010001000010010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011010001010101010101010101011001101000100110111100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111101110111011101110111011101110111011101110111011101110111111101110111011101110111011111110111011101110111011111111111111111111111111111110111011101110111111111111111011101111111111111111111111111111111111111111111111111110111011111111111111111111111111111111111111111110111111111111111111111111111111111111111011101111111011101110111111111111111111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101111011111111111111111111111111111110111011011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110011001100110011001011110010111100110010111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111100110010111100110011001100110011001101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100101110111011101110111010100110011000011101111000100110101011101110111011101110111011101110111011101110101010100110001000011101100101010000110011001100110011010101010101010101100110011110001000100110011001101010111011101110111011101110101001100110011001100110011001101010101010101010101011,
	2400'b001000010001000100010001000100010001000100010010001000110101011101111000100001010100010000110011001101000100001100100010001000100010001000100010000100100010001100110010001000110111011101000001001000100010001000100010001000100010000100010001001000100001001000100010001000100010001000100010001000100010001000100010001100110011001100110100010001000101010101010101010101010101010101100110100010101011110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011101111111011101110111011101111111011101111111011111110111111111111111111111111111011101110111011111111111011101110111111111111111111111111111011101110111111111111111011111111111111111111111111101111111011101110111111101110111011101110111111111110111011111110111011111111111011111110111111111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111011101101110111011101111011111111111111101111111111111110111011011101110111011101110111001101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011110010111011110011001100110011001101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100101110101010101010101010101010001000100001110111100010001010101110111011101110111011101110111011101110101001100110000111011001100101010000110011001100110011010101010101010101100111011101110111011110001000101010111011101110111011101010011001100010001000100110011010101010101010101010101010,
	2400'b000100010001000100010001000100010001000100010001000100010010001101000101011001010101010101000100010001000101010100110010001000110011001100110010001000100011010001010101001000100101100001000010001101000011010000110010001000100010000100010001000100100010000100100010001000100010001000100010001000100010001000100011001100110011010001000100010001000100010001000101010101010101010101010101010101010110011110011011110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011111111111011101110111011111111111011101110111011101110111011101111111011111110111111111111111111111111111011111110111011101110111011101110111011111110111111101110111011101110111111111111111111111111111111111111111111111111111111101111111111111111111111111110111011101110111011111110111111111111111111111111111111101110111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011101110111011101111011111111111011101111111111101110111011011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110010111011101111001011110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111100101110111011110011001100110011011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100101110101001100110101010101010011000100001110110011110001001101010111011101110111011101110111010101010101001100001110111011001010101010000110011001100110011010101010101010101100110011001110111011101111000100110111011101110111010100110001000100010001001100110101010101010101010101010101010,
	2400'b001000010001000100010001000100010001000100010001000100010001000100010010001000110100010101010101011001010101010000110011001100110011001100110100001100100011010101100111010000100010011000110001010101100100010100110010001100100010000100010001000100010010001000100010001000100010001000100010001000100011001100110011010001000100010001000100010001000100010001000101010101010101011001100101010101010101011001100111100010101100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101110111011111110111111111110111111111110111011101110111011101110111111101111111111101110111111111111111111111111111111111111111011111110111111111111111111101110111111101111111011101110111011111110111111111111111111101111111111111111111111111111111111111110111011111111111111111111111111101111111111111111111111111110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111011101110111011110111111111111111111111110111011101110111011011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001011110010111011110011001100110011001100110011001100110011001100110011001100110011001100101110111100101110111011101111001100101110111100110011001100110011011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110010111010100110011001100110011000100010000110011001111010101010111011101110111011101110101010100110011000011101110110011001010100010000110011001100110011010101010101010101010110011001110111011110001000100110111011101110101001100010000111100010011001100110101010101010101010101010101010,
	2400'b001000100001000100010001000100010001000100010001000100010001000100010001000100010010001000110100010101010101010000110011010101010011010001010110010101000011001101110110010100100010001100100010011001110101010000100011001100100010000100100001001000100010001000100010001000100010001000100011001100110011001101000100010001000100010001000101010101000100010001010101010101010101010101010101010101010101010101100110011101111000101010111101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111111110111011111111111111111110111011111111111111101110111011111110111011111111111111111111111111111111111111111111111111111111111111111110111111101110111111111111111011101111111011111111111011111111111011111111111111111111111111111111111111111110111011111111111011111111111111101111111111101110111011111111111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111101101110111011101110111011110111011101110111111111110111011111110111011011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001100110010111100110011001100110011001100110011001100110011001100110011001100110011001100110010111100110011001011110011001100110011001100110011001100110111011101110111011101110111011101110111001100110011001100110011001101110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110010111010101010011000100010001000011101110111011001101000100110101011101110101011101010101001100010001000011101100101010101010100010000110011001100110100011001010100010101010110011001100111100010001001101010101010101010011000011101111000100010011001100110101010101010101010101010101010,
	2400'b001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001101000100010000110011010001010110010101111000100001110101001001011000011000110001000100100010010101010100001100110011001000100001000100100001001000100010001000100010001000100010001100110011001100110100010001000100010001000100010001010101010101010101010101010101011001100110011001100101010101010101011001100110011001111000100010001001101011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101111111011101110111011101111111111111111111111101110111011101110111011101110111011101111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111101101110111011101110111011101110111011101111111111110111011101110111011011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011100110011001100110011001100110011001100110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111001100110011001100110011011100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001011101010101001100001110111100001110111011101010110100010011010101010101010101010101001011101100110011001100101010101000100010000110011001100110100010101000100010101010110011001100111011110001001101010101010100110000111011101111000100010011001100110011010101010101010101010101010,
	2400'b001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001100110100011001010110011001101000100110000111010000110111011100110001000100010010010000110010001100110010001000010001001000100010001000100010001000100010001000110011001100110011001101000100010001000100010001000101010101010101010101010110011001100110011101110111011101110110011001100101011001100110010101101000101010111010100110001001101011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011101101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111011101110111111111111111011101111111111101110111011101110111111111111111111101111111111101110111011101110111011111111111111101111111011101111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111101101110111011101110111011101110111011101111011111111111111111110111011101101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011110110111011101110111011100110011001100110011001101110111011101110011001100110011001100110010111100110011001100110011001100110011001011110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001100110011001101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101010101010100110000110011110000111011101100100011101111010101010101010101010101001100001100110010101010101010101000100001100110011001100110100010101000100010101010110011001110111011110011001101010101001100001110110011001110111100010001000100110101010101010101010101010101010,
	2400'b001000100010001000100010001000010010001000100001000100010001000100010001000100010001000100010001000100100010001000100011010001100101010101010101100010001000011000100100011101010010000100010010001100100011001100100010001000100010001000100010001000010010001000110011001100110011001100110011010001000100010001000100010001010101010101010101010101100110011101110111100010001000100110001000011101100110011001110111011001100110100010101100110010111001100010001001110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101111011011101110111011101110111011101111011101101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111011101111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111110111111101110111111111111111011101110111111111111111011101111111011111110111011101110111011101110111011101110111111111110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111110111111111111111111111110111111101101110111011101110111011101110111011101111011111110111011101110111011101101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111101110111011101101110111011100110011001100110011001101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101010101010100110010111010101100111011001100100011001111000101010101010101010101001011101100110011001010100010001000100001100110011001100110101010101000100010101010110011101110111100010011001100110011000011101100110011001100110011101111000100110011010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100100011001100110010001000110100010101110110010001111001011100110010011001100010000100010010001100100100001100100001001000100010001000100010001000100011001100110011001100110011001100110011010001000100010001000100010001010101010101010101010101100111100010001000100010011001100110011001100010001000011101110111011001100110011101111001101111011101110010101000100010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110111011011101110111011101110111011101111011101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111011101110111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111110111111111111111011111110111011111111111011101110111011101110111111101111111111111111111111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111101110111111111111111111111111111111101101110111011101110111011101110111011110111011111110111011101110111011011101111011101101110111011101110111011101110011011101110111001100110011001100110011001100110011001100110011001100110011001101111011101110111011101110111011011100110011001100110011001101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110011001100110011011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110101001100110011000011101100101011001100101010001100111100110101010101010101001100001110110010101010100001100110011001100110011001100110100010101000100010101010110011101110111100010001001100110000111011001100110010101100101011001111000100110011010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001100100010001000100010001000010001000100010001001000100010010001000100010000110010001101011000011101010111100001010010010001010010000100010010001000100101001100100010001000100010001000100010010001010101010000110011010001000100001101000100010001000100010001000100010001000101010101010101010101100110011101111000100110011001100110011001100010001000100010000111011101100110011001100111100010101100110111011100101010011001101111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011101110110111011101110111011101110111011101110111011110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111111111011101110111011111111111111101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011011101110111011101110111011101111011101110111111101110111011101110111011101110111011101101111011101101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011011101111011101110111011101110111011011101110011001100110011001100110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001100110011011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111010100110001000011101100101010101000101001101010111100010101010101010101001100001110111011001010100010000110011001100110011001100110100010101000100010101100111011001110111100010001001100001110110010101010101010101010101011001111000100010011010101010101010101010101000,
	2400'b001000100010001000110011001000100010001100110100001100110010001100100010001100110010001000100010001100110011001100110100011001110101001000100100011001110101011001010010001001000010000100010010001001000100001000010010001000100010001101000101011101100100001101000100010101000100010001000100010001000100010001000100010001000100010101010101010101010101010101100111100010011010100110011010100110001001100110011001100001110111011001110111011110001001101111011101110111001010100110101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011101110110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111101110111111111111111111111111111111111111111011111110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111001100110011001100110011001100110011001100110011001101110111011110111011101110111011101110111011101101110011001100110011001100110011011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101111001100110011011101110111011101110111011101110011001100110010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111010100110011000011101110110010101000100001100110101011110011010101010011001100010000111011001010100010000110011001100110011001100110100010101000100010101100110011001110111100010001000011101100110010101010101010001010101011001111000100110011010101010101010101010011000,
	2400'b001100100011001101000011001000110100010001100110010000110100010000110100010001000100001100100100011001010101010101100101010101100111011101000010001001000101010001000011001000110010000100010010001001000011001000010010001000100011010001010100010000110011010001010101010101010100010001000100010101000101010101000100010001000100010001010101010101010101010101010101011001100111011110011001100110011001100110011010100110011000100010001000100010001001101011001101110111011101101110011001101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011100110011001100110011001100110111011101111011101110111011101110111011101110111011011101110011001100110011001100110011011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101111001100110011001101110111011101110111011100110011001100101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101010011000100001100110010101000100001100110100011010001001101010011001011101110111011001010100010000110011001100110011001100110100010101000101010101010110011001110111100010000111011001100101010001000100010001010110011001111001100110101010101010101010100110001000,
	2400'b001100110100010101000011001101000101011110011000010001000110010101000100010101000100001100100110100001110111100010011000100110000111011101110110001100100010001100100010000100100010000100010001001001000010000100010001001000100011001100110011010001010110011101110110011001100101010001010101010101010101010101010100010101010101010101010101011001010100010001000100010101010101010101010110011001100111100010011010101010101001100110011000101010101011101110011100110111011101110111001010100110011010110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111111101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111011111111111111111111111111111111111011101111111011111111111111101111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111110110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111111101110111011101110111011101101110111011101110111011101110111011101110111001100110011001100110011001100110111011101111011101110111011101110111011101110110111011100110011001100110011001100110011001101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101111001100110011001100110111011100110011001100110011001100101110111011101111001100110011001100110011001100110011001100110011001100110011001100110010111100110011001100110011001100110011001100110011001011110011001100110011001011110011001100110011001100110011001100110011001011101010011000100001110110010101010100010000110011010101111001100110011000011001100110010101010100010000110011001100110011001100110100010101000100010101010110011001110111011101110110011001010100010001000100010101010110011110001001100110101010101010101001100010001001,
	2400'b001101000110011101010100010001010111101010100111010001110110010101010110010101010100001100100111100110001001101010111010101111001011100010001000011000110010001000100001000100010001000100010001001000100010000100010001001000100011010101100110011001111000011101110110011101110101010101010101011001100110011001010101011001100110010101100110011001100101010101010100010101010101010101010101010101010101011001101000100010011001101010101001101010111011101010001010110111011101110111011101110010101000100111001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111101101110111011101110111011101110111011101110111011101110111011101110111101110111011111111111111111111111111101110111011101110111011101110110111011101110111011101110111011101110111001100110011001100110011001100110111011101110111101110111011011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101111001100110011001100110011001100110011001100110011001011101110111011101111001100110011001100110011001100110011001100110010111011101110111100101111001100110011001100110011001011101110111011101110111011101110111011101110101010101010111011110011001100110011001100101110111010101010101001100001110111011101010100001100110011001101011000100110011001011101100100010001000100010001000011001100110011001100110100010001000101010101100110011001110111011001100110010101000100010001010101011001111000100110011010101010101010101010011000100110011001,
	2400'b010110001010100001010101010101011001101110010101011110000101011001110110011001100011001000111001100110011010101110111011101111001100101110101011101001110100001000010001000100010001000100010001000100010001000100010001000100100110100110101001011101100110011101110111011001100100010001010101011010000111011001010101011010001000011001110111100001110110011101100101010101100101010101010101010101010101010101010101010101100111100010101010100110011001100010001000101111011101110111011101110111011011100110011011111011101110111011101110111011101110111011101110111011101110111011101101110111011101111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111111101111111111111110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011011101110111011101110111011101110111011101110111011101110111011101111011101110111111111111111111111111111111111111111011101110111011101110110111101110111011011101111011011101110111011101110011001100110011001100110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110010111011101110111011101110111100110011001100110011001100110011001100110011001011101110111011101111001100110011001100110011001100110011001100110010111011101110111100110011001011101010101001100001110111011001010101011001100111011101100101011101111000100110101011101110111100110011001100101110111001100010001000100010000111011001100100001100110011001101000111100110001000100001110101010000110011001100110011001100110011001100110100010001000100010101010110011001100110011001100101010001000100010101010110011110001001100110011010101010101010101010001000100110011001,
	2400'b100010111100011001101000011010001011110010010111101010010111011101100110011001010010001001001000100010101011101110111011101110111011101110101010100101110100000100010001000100010001000100010001000100010001000100010001000100100100100010011001100001110111100001110110011001010100010101010101011010000111011001010101011110011000011010001000100110000111100001110101011110000110011001100110010101010101010101010101010101010101011001111000100010011001100010001000100111001101110111011101110111011101110110111001101111101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111111101110111011101110111011101110111011101111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101101110111011101110111011101110111011101110111011101110111011101110111101110111011101111111111111111111111111111111111111111111111111111111111101110111011101110111011101110110111011101110111011101110111001100110011011101110111011101110111001100110011011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100101110111011101110111011110011001100110011001100110011001100110011001011101110111011101110111100110011001100110011001100110011001100110011001100101110111011101110101001011101100101010101000100010001000011001100110011001100110011001101000100011001111000100110101011101111001100101110111001100001110111011101110111011001100101010000110011001000110101100010000110011110000110010000110011001100110011001100110011001100110100010001000100010101010101011001100101011001100101010101010101010101100111011110001001100110011001101010101010100010001001101010101001,
	2400'b110011001010011110101000011110111101110010001011101110011000011101010110010100110010001001011000100010101010101010011001100001110111011101010011001100100001000100010001000100010001000100010001000100010001000100010001000100010010010101010101010101000100010001000100010001000100010001010101011001110111011001100101011110101001011110011001100110011000101010010110100010010111011110000111011001100101010101010101010101010101010101010110011110001001100110011001100110101100110111011101110111101101110111011100101111001110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011011101111011101110111011011110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111111101110111111101110111111111110111111101110111011101111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110110111101101110111011101110111011101110111011101110111011101110111001100110011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110010111011101110111011101110111011110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111100110011001011101111001100101110111010100001110110010101010101011001100101010101010100010001000100001100110011001100110011010001000101011001111001101010111011101110111010100110000111011101100111011001100110010100110011001000110100011110000111010101100110010101000011001100110011001100110011001100110101010001000100010001000101010101010101011001010101010101010101011001100111011110001001100110011010101010101001100010011001101010011010,
	2400'b110010111000100110101001100111001101101110111100101110011000011001010100001100100010001000110100010001000100001100110010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001100110011001101000100010101010110011001100101011010011001011110011010101110111001101010110111100110100111011110000111011101110110011001010101010101010101010101010101011001111000100110011001101010101100110111101110111011101110111011011101110111011101111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011110110111001100111011101110111011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110110111011101110111011101110111011101110111011101110111011101110111011110111011101110111111111110111011111111111111101111111111111111111111111110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110011001100110011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100101110101000011101100110010101100110011001100101010101000100010001000100001100110011001100110011001100110011001101000101011010001010101110111010100110001000011101100110011001010110010101000011001100110011011010000110010101000101010101000011001100110011001100110011001101000101010001000100010001000100010101010101010101010101010101010101010101100111011110001001100110101010101010011000100110101010101010101010,
	2400'b110010101011101110101010101011011100101111001010101001110101010100110011001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000110011001100110100010001000100010001010101010101100111011010011010101110111010101110111001101010111000011101111000011101110111011101110110011001010101010101010101011001100110100010011010101010111100110111011110111011101110111011101101110111101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110110010111100110111101110111011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111111101110111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110110111011101110111011101110111011101110111011101110111011101110111011110111011101110111111101110111111111111111111111110111011111111111111111111111111101110111011101110111011101110111011101110111011011101111011011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110001000100001100111011001110110011001100101010101000100010000110011001100110011001100110011001100110011001100110011001101000101011110101011101010011000011101100110011001100110011001010100001100110010010101110110010001000100010001000100001100110011001100100010001101000101010001000100010001000100010001010101010101010100010001010101010101100111100010001001100110011001100101111000100110101010101010101010,
	2400'b101010101011101111001011110011001010101010011000011001000011001000100001000100010001000100010001000100100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100011001100110011010001000100010001000100010001000100010101101000101010111011101110111010101110111010101010011001100001110111100010000111011101110110010101010101011001100110011001111001101110111100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101011001101101110111011110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111011111111111111111111111111101111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110110111011101110111011101110111011101110111011101110111011101110111011110111011101110111111101110111011111111111111111111111011111111111111111111111111101110111011111110111011101110111011101110111011101110111011101101111011011101110111011101110111001100110111001100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001011110001000100001110110011001100101010101010100010001000011001100110011001100110011001100110011001100110011001100110011010001000110100110101001100001110110011001010110011001100101010000110010010001100101010000110011001100110011001100110011001100100010001000110100010001000100010001000100010001010101010101000100010001010101011001100111100010001001100110011001011110001001101010101010101010101010,
	2400'b101110111011110011001011101010101000010101000011001000100001000100010001000100010001000100010001000100010010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000110011001100110011001100110011010001000100010001000100010001000011001101000100010101111000101010111011110010111010101110101010101010011000100010011001100010001000011101100110010101010110011001100111100110111100110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111101110110111011101110111011101110111001100110011001100110111011101110111011101110111011101110111011101110010111001100111001100101010101011110011101110111011101110111011011100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111110111011101101110111011101110111011101110111011101110111011101110111011101110111101110111011111110111111101110111011111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011011101111011011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001101010101000100110011001100001110111011001100110011001100110010101000100010101010100010001000011001100110011001100110011001100110011001100110011010010001010101010000111011001010101010101100101010000110010001101010101010001000011001100110011001100110011001100110010001000110011010001000100010001000100010001000100010001000100010001010101011001110111100010011001100110010111011110011010101010101010101010101010,
	2400'b101110111100110010101000010101000011001000100001000100010001000100010001001000010001000100010001000100010010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100011001100110011001100110011001100110011001100110100010001000100001100110011010001000101011001111001101010111011110010111010101110101000100010011010100110011001100110000111011001010101011001100111011110101100110111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011110110111011101110111011101110111001100110010111010101111001101110111011101110111011101110111011100101110011001100110111011101010101011110111101110111011111110110010111010101111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111110111011101101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011011101111011101101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101111001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010011001100110101010100110001000100001110111100010000111010101010110011001100110011001100110010101000011001100110010001000100010001000100010001000110110100110011000011001010101010101100101010100110010001101010101010000110011001100110011001100110011001100100010001000110011001101000100010001000100010001000100010001000100010001010110011001111000100010001001100101110110100010101010101010101010101010101010,
	2400'b101110011000011001000011001000100001001000010001000100010001000100010010001000010001000100010001000100100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100100010101000011001100110011001000100010001100110011001100110100010001000100010000110011001100110100010001000011001101000100010001010110011110001001101111001011110010111001100110011010101010101010101110101000100101110110010101100110011001111011110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110011001100101110101010101010111100110111011101110111011101110111001011100110001000100010101010101010101011110011101110111011011011101010101010101111011110111011101110111111101110111011101110111011101110111011101110111011111111111011101111111011101110111011101110111111111110111011111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011110110111011110111011101110111011111111111111111111111111111111111111111111111111111111111111101110111111111110111011101110111011101110111011101110111011101110111011011101110111001100110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101111001100110011001100110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001101010111011100110011010100110011001101010010111011110001000100010001000100010000111011001010100001100110011001000100010001000100010001000100010010110001000011101110101010101010101010001000010001001000100010000110011001100110011001100100011001100110010001000110011001100110100010001000100010001000100010001000100010101010110011001111000100010001001100001100111100110101010101010101010101010011001,
	2400'b011001000010001000100010001000100001000100010001001000010001000100010010001000100010000100100001001000100010001000110010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010010001000100100011001100110010101000011001100110011001100110010001100110011010001000100010001000100010000110011001100110011001100110011010001000101011001100111100010011010101111001011101010011010101110101010101110111001101010010111011001010110010101100111101111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011100110011001011101110101010100110011011110111011101110111011101110111001010100110001000100010011001101010101011110111101110110110111010101010101010101111011110111011101110111111101110111111111110111011101110111011111111111011101110111111111110111011101110111011101110111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101111011101110111011101110111011101111111111101111111111111111111111111111111111111111111111111111111111101111111111111111111011101110111011101110111011101110111011101101110111001011101110111011101111001101110111011100110011001100110011001100110011001100110011001100110011001100110011001100101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101111001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111011100110111011101110101011101110111010101010101010101010101001100010000111011101010101010000110011001000100010001000100010001000100010001000110110100001110110010101010101010001000010001001000101001100110011001100110011001100100010001000100010001100110011001100110011010001000011001101000100010001000100010101010110011101110111100010000111011001111000100110101010101110111010100010001010,
	2400'b001000100010001000100010001000010001000100010001001000100001001000100010001000100010001000100001001000100010001000100010001000100010001000100001000100010010001000100010001000100010000100010001000100010001001000100011001000110011010101101000100001110110010101000100010000110011001100110011010001010110011001010101010101000011001100110011010001000011010001000101010101010110011101111000100010101010101110111010110011001011101111001010101110111001011101100110011001010101100011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110011001100110011001011101110101010100110011010101111011101110111011101110111001001100010001000100010011001100110101100110111101101101110101010101010101010101111001110111011101110111011111110111011101111111011111110111011111111111011101110111011101110111011101110111011101110111111111110111111101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011111111111111101110111011101110111011101110111011011101110111011101110111011101110111101101111011101110111011101110111011101110111011101110111011101110111111111111111011111111111111111110111011111111111111111110111111101110111011101110111011101110111011101110111011011100110011001011101010111011101110111011110111011100110011001100110011001100110011001100110011001100110011001100110011001100101110111011110011001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101111001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111100110010111100110011001011101110111011101110011000100001110110011001010100010000110011001000100010001000100010001000100010001000100010010001100110011001010101010001000010001000110101001100100011001100110011001100100011001000100010001100110011001100110011010000110011001101000100010001000100010101100110011101110111100010000110011010001001101010101011100101100110100110101010,
	2400'b001000100010001000100010001000100001000100010010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100100010001000100010001000100010000100010001000100100010001001000100001100110100001101000110100010011000100001110101010101010100010001000100010101100111011101110110011001010100010001000100010001000100010001000100010101010110011001110111011110001000100110101010101111001100101111001011101111001011100101110111011101100101011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110011001100110011001011101110111010100110011001101010111101110111011101110111001010100010001000100010011001100110101100111011011010101010101010101010101011110011011110111011101110111111111110111011101110111111111110111011101110111011101110111011101110111111101110111011101110111011111110111111101110111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111101110111011101110111011111111111011101110111011101110111011101110111011101101110111011101111011011110110111101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111111110111011111110111111111110111011101110111011101110111011101110111011101110110111011100110010111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111010101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100101111001011101010000101010101010101010101010100010000110011001000100011001000100010001000100010001000010001000100100100011001010101010101000010001000110101010000110010001000110011001100100010001000100010001101000100001100110011010000110011001100110100010001000100010101100110011101111000100001110110100010011010101010010110010001101001101010011001,
	2400'b001000100010001000100010001000100010001000010010000100010010001000100010001000100010001000100010001000110011001000110010001000100010001000100010001000100010001000100010001000100010001000100010000100100010001001000101010100110011001100110100011001111001101010101001011001101000011001100110011001100111011101110111011001100101010101000100010001000101010101010100010001010110011001110111011110001000100110011001100110111100101111001100101011001011101110000111100001110101010101111100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011100110010111011101110111011101110111011101010011000100110101100110111011101110111001001100010001000100010011001101010111101110010101010101010101010101010111100110011011110111011101110111011111111111011101110111111111111111011111110111011101110111011101110111011101110111011101111111111111111111011101110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011111111111111101110111011101110111011101110111011101110111011101110111011101110111011011110110111011101111011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101110111011101110111011101110111011101110110111011100110011001100110011001100101110101010100110101011110011001100110011001100110011001100110011001100110011001100110011001100101110101011101110011010101110101011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100101110111011100110000111011001100101011001010101010000110011001101000100001100100010001000100010001000100010000100010010010001010101010101000011001000100100001100110010001000100010001100110010001000100010001101000100001100110011001100110011001100110011010001000100010101100110011001110111011101100111100010101010011101000100100010101010101010010111,
	2400'b000100010010000100010001001000100010001000100010000100100010001000100011001100100010001000100010001101000011001100100010001000010001001000100010001000100010001000100010001000100010001000100010001000100010001000100100010101010011001100100011010001010111100110101011101010001000100110000111011101110111100010001000011101100101010101000101010001000101010101010101010101010101011001110111011101111000100010011001100110011010101111001100101111001100101110111000011110000110010101100111110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111001100101110101010101010101010101110111011101110101001100010011010110011011101110111001010100010001000011110001001101011001100101010011001101010101010101111001101110111101110111011101110111011111110111011111111111111101111111111111111111111101111111111101110111011111111111011111111111111101110111011101110111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101101110111011101110111001100110011001011100110000111011001111000101011001100110011001100110011001100110011001100110011001100110011001100101010101010101010001001100110011001101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100101110111001100010001000011101110110010101010100010001000101010101000011001100110010001000100010000100010001000100010001000100110100010101000011001000100010001100100010001000100010001000100010001000100010001101010101001100100011001100110011001100110011010001000101010101100110011101110110010101101000100110010101001101011001101010101010100101110101,
	2400'b000100010001000100010001001000100010001000100010001000100010001100110011001100110011001000100011010001000100001100100010000100010001001000100010001000100010001000100010001000100010001000100010001000100010000100010011010101100100001100110010001101000101011010001011110010111000100010011000011110000111100010001000100001110110010101010101011001000100010001010101010101010110011001100111011110001000100010001001100110011010101111001100101111001100110011001010011110000111010101100101011111001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111001100101110101001100110011001100110011001101010111010100110001001101011001101110111001010100001110111011110001001101010111010100110011010101010101011110011011110111011101110111011101110111011101110111111101111111111111111111111111111111111111111111111101110111011111110111011111111111111101110111011101110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111001100110010111001100001100101010101010101011110101100110010111011110011001100110011001100110011001100110011001011100110011001100010001001100010001001101010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011101110011000100010001000100001110111011001100101010101100101010001000100001100100010001000100001000100010001000100010001000100010010001101000011001000010001001000100010001000100010001000100010001000100010001101000101001100100011001100110011001100110011010001000101010101100110011101100101011010001001011100110100011110011001100110101001011001010100,
	2400'b000100010001000100010010001000100010001000100010001000100010001100110011001100110011001000110011010000110011001000100010000100010010001000100010001000010001000100100010001000100010001000100010001000100010000100010011010001010101010000110011001100110101011001100111101010111011011101111000100110011000100010011001100110000110011001010110011101010100010001000101010101100110011001100110011101111000100010001000100010001001101010111100110011001100110011001011100010000111011001100110010101111100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100101110111010100110011001100110001000100010001001100110011001100110101101110111001001100010000111011101111000100110001000100010011001100110101011110111101110111011101110111011101110111111111110111111111111111111101110111111111111111111101111111111101111111011101110111111101110111011101110111011101111111111101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110111011110111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011111110111011111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110010111001011101100101010101000100010001101010101110011011110011001011110011001100110011001100101110101001100010000111011110001000100010001000100110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011101010011000100010001000011101110111011001010110011101100101010001000100001100110010001000100001000100010001000100010001000100010001001000100010000100010001001000100010001000100010001000100010001000100010001101000100001100100010001100110011001100110100010001000101010101010110011001010101100010010110001101011000100110101001100010000111011001010100,
	2400'b001000010001000100100010001000100010001000110010001000100011001101000100010001000100001100110100010000110010000100010010001000100010001000100010001000010001000100100010001000010001000100100010001000010001000100100011010001000101010101000011001100110011010101100110011001111001100110001000100010011000100010011001100110001000011101100110100001100101010001000101010101010110011001100110011001100111100010001000100010001000100110011011110011011100110011001100101010000111011001100111011001011000110011101101111011101110110111011110111011101110111011101110111011101110111011011101111011101110111011011101110111011100110011001100101110111011101110101001100110011001100001110111011110001001100110011011110011001010100010000111011101111001100110001000100010001000100110101100111011101110111011101110111011101110111011101110111111111110111111111111111111101110111011101110111011111111111111111110111011101110111011111111111011111110111011101110111011101111111111111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110111011100110011001100110111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011111111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011100101010011000100001110110010101000100010001010111101010001000101110111010101111001100110011001011100101110111011001110110011001110111011101111001101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011000100010001000100001110110011001110110011001100110010101000100001100100011001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001101000011001000100010001100110011001100110100010001000100010101010101010001011000100101010011011010011010101010011000011001110101010101000100,
	2400'b001000100001001000100010001100100010001000110011001000110011010001000100010001000100001100110100010000100010000100100010001000100010001000100010001000010001000100100010001000010001000100100010000100010001000100100100011001010101011001010100001100110011001101010111100001100101011101111000100010001000100010001001100110011000100001110111100110000110010101010101010101010101011001100110011101110111011110001000100110011000100010011010110011001100110011001100101110101000011001110111100001100101100111011101110111011101110111011110111011101110111011101110111011101110111011101101110111011101110111011101110111001100110011001100110011001011101110111001100110011001100010000111011001100111100110011001101010111010100001110111011101111000100110011001100010001000100110111100110011001101111011101110111011101110111011101111111111111111111011111110111111101110111011101110111011101110111011101110111111101110111111111110111011101110110111011110111011101110111011111111111111111111111111101111111111111110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110011001100110011001100110011001101111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110110111101110111011101110111011101110111011101110111011101110111011101101110111001011101010101001100001110110010101010100010001000101100010000110100010101001101010111011101110111001011101100101010101100110011001100110011110001010110011001101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111010100110001000100010001000100001110111100001110111011101110110010101000100001100110011001000100010000100010001000100010001000100010001000100010001000100010001000100010001001000100001000100010010001000100010001101000011001000100011001100110011001100110100010101010101010101010100010101111001011001001000100110011001100001100101010001000100001100110011,
	2400'b001000100010001000100010001100110011001001000011001100110100010001000101010001000100001100110100001100100001000100100010001000100010001000100010001000010001000100010010001000010001000100010001000100010001000100100101011101110101011001100101010000110011001101000110011101110110010101010110011101111000100010001001100110011001100010001000101010010111010101100101010101010101010101010110011001110111011110001000100010011001100110011001101011001101110111011100110010111001011110001000100010000110011010011100110111011101110111011101111011101110111011101110111011101110111011101101110111011101110111011101110111001100110011001100110011001100101110111010100110011001100110000111011001100110011110011000100010101001100001100110011001100111011110001000011110001000100110101010100110011010101111001101111011101110111011101111111111101111111011111111111111101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101111011101110111011101110111111111111111011101111111011101110110111101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011100110011001100110011001100110011001100110011001101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111101110111011101110111011101110111011101110111011011101110111011100101110111010100001110110010101010100010001000100011001100101011010001000100110101011101110101000011001010101010101010101011001100111100010101011110011001100110111011100110011001100110011001100110010111100110011001100110011001100110011001100110011001100110011001011101110111011110010111011101111001011101111001100101110111011101110111011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110001001100110011001100010001000100001111000100001110111011001010100001101000011001000100010000100010001000100010001000100010001000100010001000100010001000100010001001000100001000100010001000100010010001000110011001000100010001100110011001100110100010101010101010001000101011110000111011010001001100110000110001100110011001000100011001100110011,
	2400'b001000100010001000100010001100110011001001000100001100110100010101010101010101000101010000110011001000010001001000010010001000100010001000100010001000010001000100010010001000100010001000010010001000100001000100100110100010010111011001110111010101000011001100110100011001111000011101100110010101010110011110001001100110011001100110011000100110101000011001100110011001100110010101010101010101100110011110001000100110011001100110101010101010111101110111011100110010111010100110011010100110000111011001111010110011011101110111011101110111011101111011101110111011101110111011101110111011011101110111011101110111001100110011001100110111011100110011001011101110101001100110001000011001100110011001111000100010001000011101100110011001100110011001110111100010001000100010001000100010001001101010011010101111001110111011101110111011101111111111111111111111111110111011101110111011101110111011101111111011101110111011011101110111011101110111011101110111101110111011101110111011111110111111111110111011011101110111011101110111011110111011111111111111111111111111111111111111111111111111111111111111111111111111101101110011001100101110111011101110111011101110111100110011001100110111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111011101111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110110111101110111011101110111011101110111011011101110111011100101110101001100001110110011001010101010001000100010001010100010001100111011110001010101010010111010101010100010001010101010101100111100010011010110011001100110011001100110011001100110010111011101110101011110011001100110011001100110011001100110011001100110010111011101110111011101111001100101111001011101110111011101110111011101110111011110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011110010111001100110011001100110101010100110011000100010001000011101111000011101010100010001000011001100100010001000100010000100010001000100010001000100010001000100010001000100010001000100100010001000010001001000100010001000100010001000100010001100110011001100110100010001010100001101011000100101110111100110011000011101010011001000100010001000100011001100110011,
	2400'b001000100010001000100010001101000100001001000100010000110100010101100110011001000101010000110010001000010010000100010010001000100010001000100010001000010001000100010010001000100010001000100010001000100010001000110110100010011001011001111000011101010100001100110011010001101000100010000111011001100101010101101000100110011001101010101001100110101001011001110110011101100101010101010101010101010110011110001001100110011010101010101010101110111100110111011101110111001011101110101010101110010111011101111000101111011101110111011101110111011101110111011101111011101110111011101110111011101101110111011101110111011101110111011101110111011101110011001100110011001011101010101001100001100110010101100110011101110110010101010101010101100110011001110111011101111000100010011000100110001000100110011001100110101011110111101110111011101111111111111111111111111111111011101110111011101110111011101110111011101110111011011101110111011100110011001100110111011110111011101110111011101110111111101101110111011101110111011101110111011101110111101111111111111111111111111111111111111111111111111111111111111111111011011101110011001011101110111011101110111011101110111011101111001100110011001101111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111001100101110111010100101110101010101010101010101000011010001000100010001000101010101111001101010000111010101000100010001010101011001100111100010011010110011001101110111001100110011001011101110101001100110101011110011001100110011001100110011001100110011001100110010111011101010111011101111001100101110111100110010111011101111001100110011001100110011001100101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010111011101110101001100110011000100010011000011001010101010101000100001100100010001000100010000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100011001100110010001000100010001000110011001000100011001100110011010001111000100010001001100110000110001100100010001000100010001000100010001000110011,
	2400'b001000100011001100110010010001000100001101000101010000110101011001100110011001010100010000100010000100100001000100010010001000100010001000100010001000100001000100010001001000100010001000100010001000010001001000110101011110011010100101111000100101110100001100110011001101001000100110011001011101100110010101010110011110011010101010101010101010111010011110000111011101100101010101100101010101010101011001111000100110101010101010111011101110111011110011001101110111011100110111001011110010111000100010101000100111001101110111011101110111011101110111011101110111011101110111101110111011101110110111011101110111011101110111011101110111011101110011001100110011001100101110111011101001110101010101010110011110000110010101010101010101010110011001100111011110001000100110011010100110001000100110011001100110101010110011101110111011101110111011101110111111111110111011101110111011101110111011101110110111011101110111011101110111001100110011001100110011011110111011101110111011101110111011101101110111001101110111011101110111011101110111101110111111111111111111111111111111111111111111111111111111111110111011001100110010111011101110111011101110111011101110111011101110111011110011001100111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110111111101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011011101110010111011101010010111010101000100010001000100010000110100001101000100010101101000100110000110011001000100010001000101010101100111100110101011101111001100110111001100110010111010100110001000100110101011110011001100110011001100110011001100110010111011101110111011101110111011101110111011110011001100110010111011101111001011110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111010101010101011101111001100110010111010101010011001100110011000011101100111011001010100001100110100010000100001000100100001000100010001000100010001000100010001000100010001000100010010001000100001000100100011010001000011001000100010001000100010001000100011001100110100011110000111011110001000011001000010001000100010001000100010001000100010001000110011,
	2400'b001100110100010001000011010001010100001101000101010101000110011001100111011001000101001100100010000100010001000100100010001000100010001000100010001000100001000100010001000100010001000100010001000100010001000100110110011110001010101010010111100010000101010000110011001000110101100010101010100001100111011101100101010101111001101010101010101110111010011110010111011110000110010101100101010101010101010101100111100010101010101010111011101110111100110011001101110111011101110111011011110111001011100010111011100110011100110111011101110111011101110111011101110111011101110111011110111011101110111011011101110111011101110111011101110011001100101110111011101110111011101110101011101110100111010101010110011001111000011001010101010101010110011001110111011101110111011110001001100110001000100010011001100110011010101111011110111011101110111011101110111111101110111011101110111011101110111011101101110011011101110111011101110011001100110011001100110011011101111011101110111011111110111011011101110011001101110111011101110111011101110111101110111011111111111111111111111111111111111111111111111111111110110111001100110010111011101110111011101110111011101110111011101110111011101110111100110111101111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111111101111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111101110111011101110111011101110111011101110111011101110111011011101110111011101110011001011101010101001011001000011001101000100001100110011001100110100010001010111011101110110010001000100010001000101011001100111100110101011101110111100110011001100101010011000011101110111100110101011101111001100110011001100110011001100101110111011101111001011110011001100101110111100110011001100110011001011110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111010101110111011110011001100110011001100101010101010101010011000100010001000011101100100010001010110010100110010001000100001000100010001000100010001000100010001000100010001000100010001000100100001000100010010001000110010001000100010001000100010001000110011001101000110011101110110010101010011001000100010001000100010001000100010001000100010001000110011,
	2400'b001100110100010101010100010001100110010001000100010101000110011101110110010101010100001100100001000100010010001000100010001000100010001000100010001000100001000100010001000100010001000100010001000100010001000100110110011010001001101010101010100001110110010000110011001100110011011010011010100110000110011101110110010101100111100110101011101110111011100010011000100010000111011001100101010101000101010101010110011110011001101010101011101111001100110011011101110111011101110111011100110111011101101010101100101110011010110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001011101110111011101110101010100110011001101010101001011001010101010101100111011001010101010101010110011001100110011001100111011101111000100110011000100110011010101010101010101111001110111011101110111011101110111011101110111011101110111011101110111011101101110011001101110111001100110011001100110011001100110011001101110111101110111011101110110111011101110111001101110111011101110111011101110111101110111111111110111111111111111111111111111111111111111111101110110111001100101110111011101110111011101110111011101110111011101110111011101110111100110011011110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011001011101110101010101010101011110011011110111011101110111011101110111011101110111011011101110111011101110011001100101110111001100001100100001100110100001100110011001100110011010001000101011001110110010001000100010001000101010101100111100010011010101010101011110010111010100001110110011001100111100010011011110011001100110011001100110010111011101110111011101111001011101110111100101110111011101111001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101111001011101111001100110011001100110011001100110010111011101010001000100010011000100001100101011110000111010100110011001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001100110011010001010110010101000011001000100001001000010010001000100010001000100010001000100010001000110011,
	2400'b010001000100010101010101010101110110010101000101011001010110011101100101011001010100001000010001000100010001001000100010001000100010001000100010001000100001000100010001000100010010000100010001000100010001000100110110011110001000100110101011101001110101010001000011001100110011010001101001100110011000011001111000011101100110011110011010101111001011100110101000100010001000011001100110010101000100010101010101011010001001100110101011101111001100110011011101110111011101110111011101110111011101110010111100110011001010100110111101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110010111011101110111011101010101001100110001000100010001010100001100101010101100110011101010101010101010110011001100110011001100110011001111000100010011001100110011010101010101011101110111101111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001100110011001100110111011101111011101101110111011101110111011101110111011101110111011101111011101111111111111111111111111111111111111111111111111111111111101110110010111011101110111011101110111011101110101011101110111011101110111011101110111011110011001101111011111111111111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110111111101111111011101110111011101111111011101110111011101110111011101110111011101110111011101101101110101001100110011000100010001000100110101011110111101110111011101110111011101110111011101101110111011100110011001100101110101001100001110110010000110011001100110011001100110011010001000100010101100101010001000101010101000101010101100111100010011010101010101011101110101000011101110111011001100111100010101011101111001100110011001100101110111011101110111011101110101010101010101010101010101010101110111011101111001100110011001100110011001100110011001100101110111100110011001011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100101110101001100110101001011101111000100001110110010101010011001000100011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001100110011010101010011001000100001000100010001000100100010000100010010001000100010001000100010001100110011,
	2400'b010001000100010101010101010101110111010101000110011001010111011001100110011001010011001000010001000100100010001000100010001000100010001000100010001000100010001000010001000100100011001000010001000100010001001000110110011110001000100110101011101010010110010001000011001100110011001101000111100110011001011101101000100101110110011001111001101010111011101110111000100010011000011101110110010101010100010001010101010101101000100110011010101010111100110011011101110111011101110111011101110111011101110111011101110111011100101010011011110111011101110111011101110111011100110111001100110011001100110011001100110011001100110011001100101110111011101110111011101010011000100001110111011101110111100010000110010101010110011001010101010101010101011001100110011001100110011101111000100110011001100110101010101110111011101111001101111011101110111011101110111011101110111011101110111011101110111011011100110011001100110011001100110011011101110111001100110011001100110011001101110111011101110111001101110111011101110111011101111011101110111011101111111111111111111111111111111111111111111111101110111011101101110010111011101110111011101110111010101010101010101010111011101110111011101110111011101111001100110111101111111111101110111011101111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011011011101010011001100010001000011101110111011110001000101011001101111011101110111011101110111011101110110111011100110111001100101110101010100110000111010101000011010000110011001100110011010001000100010101010100010001000100010101010101010101100110011110011001100110101010101010000111011001100110011001100111100010101011110011001100110011001011101110111010101010101001100010000111011101111000100110011010101010101011101111001100110011001100110011001100110011001100110010111100101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110010111011101110111000100010011001100001110110011101010100001101000011001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100011001100100010000100010001000100010001000100010010001000100010001000100010001000100010001100110011,
	2400'b010001010101010101100110011001111000011001010111011101100110011001110110010101000011001000010001000100100010001000100010001000100010001000100010001000010010001000100001001000100011001100100001000100010001001000110110011110001000100110101011101010101000010101000100001100110011001100110100011110011001100101110110100010000110011001100111100010011010101111001010100110101000100010000110011001010101010001010101010101010110100110101010101010111011110011011101110111011101110111011101110111011101110111011101110111011101110110111001101011011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111010100110001000100001110111011101110110011001110110010101010101010101010101010101010101010101010110011001100111100010001000101010101011101110111011101111001100110011001101111011101110111011101110111011101110111011101110111011101110111011001100110011001101110111001100110011001101110011001100110011001100110011001100110011011101110111011101110111011110111011101110111011101110111111111111111111111111111111111111111111111111111111101110111011101101101110111011101110111011101110101010101010101010101010101011101110111011101110111011101110111100110111101111111111101110111011101111111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001100101110101010100110011001100010001000100010001001101111011110111011101110111011101110110111011101110011001100101110011000011101110111011001010100001101000011001100110011010001000100010101010100001100110100010001010101010101010110011110001001100110011001100001110110011101100101011001100110100010101011110011001100101110111011101110101001100001110111011101110111011110001001100110101011101110111011110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100101110111100110011001100110011001100110010101001100110011001100001110111011001010101010001000011001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100001000100010001000100010001000100010001000100100010001000100010001000100011001100110011,
	2400'b010101010101011001100110011110001000011101011000011101100110011101100110010101000011001000010001000100100010001000100010001000100010001000100010001000010001001000100001000100100010001100100001000100010001001000110110011110001000100110111011101010011000011000110100001100110011001100110011010010001010100110010110011110011000011001010110011101111001101111001100101010101001100010010111011101100101010001010101010101010101011110101100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011100100110101101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110101010100110011001100010001000100010000111011001010101010101010101010101010101010101010101010101100110011001111000100001111000101010111100110011001101110011011101110111011110111011101110111011011101110111011110111011101110111011101110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111101110111011101110111011101111111111111110111111111111111111101111111011111111111111101110111011101100101110111011101110111011101010101010101010101010101010101010101110111011101110111011101110111011110011011110111011101110111011111110111011101110111111101111111111111111111111101101110111011110111111111110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110010111010100110001000011101110111011101100110011110001010110011101110111011101110111011011100110010111011101010101001100001110111011001010100001100110100001100110011010000110100010001000011001100110100010001000101010001010110011110001000100010011000100001110111011001010101011001100111100110111100110011001011101110111010100110000111011101100111011001100110011101111000100110101010101110111100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001011101110111011101110111011110011001100110010111010100110000111011101100101011001100101010000110011001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100001000100010001000100010001000100010001000100010010001000100010001000100011001100110011,
	2400'b010101010110011001100110011110001000011101101000011101100110011001100101010101000010000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010000100010001001000110110100010001000101010111010100110000111011001000011001100110011001100110011001101011000101010101000011110001001100001100110011001111000100010111100101110111001100110011000011101110110010001000101010101010101011001111011110011011101110111011101110111101101110111011101110111011101110111011101110111011101110111011101110010011100110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101010101010101010101001100110011001100001110111011001010101010101010101010101010101010101010101011001100110011101111000100010001000101010111101110111101110111011101110111011101110111011101110111011101101110111011101111011101110111011101110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101111011101110111011101110111011101110111011111111111011111111111111111111111111101110111011101110111011011100101110111011101110111010101010101010101010101010101010101011101110111011101110111011101110111011110011001101110111011110111011101110111011101110111011111111111011101101111011011100110011001100110111101101110011001101111011111111111111111111111111111111111111111111111111111111111111111111111011101111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100101110101001100010000111011101110111011101110111100010111101111011101110111011011101110010111010101010011000100001110101010101010100001100110011010000110011001100110011001100110011001100110100010000110100010001000101011001110111100001110111011101110110011001010101011001111000101010111100101110111011101010011000011001100110011001100111011101111000100010011010101010111011101111001100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011101110111010100110000111011101110110011001010101010000110011001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000010001000100010001001000100001000100010001000100010010001000100011001100110011001101000100,
	2400'b011001100110011101110111011110001000011001101000011101100110011001100101010000110001000100010001001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000010010001001000111100010001001101010101010100110000111011001010100001100110011001100110011001100110101100010101010011110001001100010000110011001100110011110011100110011001010100110101001011101110110010101010101010101010101011001101000110011011101110111101110111011101110110111011101110111011101110111011101110111011101110111011101110110101100110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111010101010101001100010000111011001100101010101010101010101010101010101010101010101100110011001100111100010001000100110101101111011101110111011101110111011101110111011101110111011101110111011011110111011101110111011101110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101111011101110111011101110111011101111111011111110111111111110111111111110111011101110111011101110111011011100101110111011101010101010101010101010101010101010101010101010101110111011101110111011101110111011101111001100110011011101111011101110111011101110111011101110110111001100110011001100110011001100110011001100110011001100110111101111111111111111111111111111111111111111111111111111111111111110111111101111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110010111011101010011000100001110111011110001000100010001010110011101110111011101110110110111010101010101001100001110110010001000011001100110011001100110011001100110011010000110011001100110011001100110011010001000101011001100111011001100110011001100110010101010110011110001000101010111011101110111001100001100110011001100111011110001000100010011010101010111011110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011000100010000111011001010100010001000011001100110011001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100100010001100110011001000100010000100010001000100010001000100100010001000100010001000010010001000100010001100110011001100110100,
	2400'b011001110111011101110111100010001001011001111000011101100110011001010100001000010001000100010001001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000100010001001011000100110011001101010101010100110000111011001010101001100110011001100110011001100110011010110001010100101111001100110010111011101100111011110001010110011001100101010101010100110000111010101010101010101010101011001100111101011011101111011101110111011101110111011011101110111011101110111011101110111011101110111011101101110111101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111010101010101001100110000111011001100101010101010101010101010101010101010101010101010101010101010101011001100111011110011100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111101110111011101110111011101110111011101110111011101111111011101101110111101110111011101110111011011011101110111010101010101010101010101010101010101010101010111011101110111100110011001011101110111011101110111100110011011101110111011110111011101110111011011100101110111011101110111011101111001100110011001100110011001100110011011110111111111111111111111111111111111111111111111111111111101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001100101110101001100001110111011001100110011110001000100010101100111011101110110110111010101010011001100101110111011001000011001100100010001100110011001100110011010000110011001100110011001100110011010001000101011001100110010101010110011001010101010101111000100001110111100110101010100101110110011001100110011001111000100010011001100110101011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010011001100110000111011001010101010001000101001100110011001100100001000100010001000100010001000100010001000100010001000100010001000100010001001000100100010001000100001100110010001000100010000100010010000100010010001000100010001000100010001000100011001100110011010001000100,
	2400'b011001110111100010000111100010011001011001111000011101010101010101000010000100100001000100010010001000100010001000100010001000100010001000100010001100110010001000100011001100100011001000100010001000100011001101011000100110011010101010101010100101110111011001100101010000110011001100110011001100110011001101011001101010001000100110011001011101110111011110001001101111001100101110111011101010011000011001010101010101010101010101100110100011001101111011101110111011101110111011101110110111011101110111011101110111011101110111011100101111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100101110111100110011001100101110101010101010011001100101110111011001100101010101010101010101010101010001000100010101010101010101010101010101100110011001111010110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111101110111011101110111011101111111111101111111011101111111011001100101111001101111011101110110111001011101110101010101010101010101010101010101010101010101111001100110011011101110111011100101110111011101110111011110011011101110111011110111011101110110111001011101110111011101110111011101110111011101111001011101110111100110011011110111111111111111111111111111111111111111111111111111111101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100101110111010100110011000100001110110011001100111011101111001110011011101110111001100101010011000011101100110010101000100001100100010001000110011001100110011010000110011001100110100010000110011001101000101010101100101010101010101010101010110011110001000100001111000101010010111010101010101010101010110011001111000100010011010101010111011110011001100110111011100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010100110000111011001100101011001100101001100110011001000100001000100010001000100010001000100010001000100010001000100010001000100010001001001000110011001100101010000110001001000100001000100010010001000100010001000100011001100110011001100110011001100110011010001000100,
	2400'b011010000111100010001000100010011000011010001000011001010101010000110001000100010001000100010001001000100010001100100010001100110011001000100010001100110010001000100010001100110011001100100010001000100100011001111000100110101010101010101010100101110111011101100110010001000011001100110011001100110011001100110101100110101000101010001001100001110111011101111000100110111100110011001011101110101001011101100101010101010101010101100110011110111101111011101110111011101110111011101110110111011101110111011101110111011101110111001100110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101010101001011101100110011001110101010101010101010101010100010001000100010101010110010101010101010101010110011001111000101011001101110111011101111011101110111011101110111011101110111011101110111011101110111011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111101110111011101110111011101110111011101111111011101110110111001011101110111011110011011101110111001011101110101010101010101010101010101010101010111011110011011101111011101110110111001011101110111011101110111011110011001101110111011101111011101110110010111011101110111011101110111011101110111011101110111011101110111100110011011110111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100101110111011101010101010100110000111011101100110011001110111100010101100110111011100101110101001011101100100010000110011001100100010001000100010001100110011001100110011001100110100010001000011001101000101010101010100010001010101010101010111011101111000100010011001100001100101010001000101010101010101011001100111100010011010101010111100110011011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010100010001000011101100110011001100101010101000011001000010001000100010001000100010001000100010001000100010001000100010001000100010010001101010110011001100101001100100001000100010001000100010001001000100010001000110011010001000100010001000100010001000100010001000100,
	2400'b011110001000100010001000100010010111011010001000011001010100001100010001000100010001000100010001001000100010001100110010001100110011001100100010001100110010001000100010001000110100001100110011001100110100100010011001101010101010101010101001100001110111011001110111010001010011001100110011001100110011001100110011011010101010101010101001101010011000011101111000100010101100110111001100110011001010011101110110011001010101010101100110100010101101111011101110111011101110111011101110111011101101110111011101110011001101110111001101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101010101000011001100111100010000110010101010101010101010100010001000100010001100111011101110110011001100110011001100111100110111100110011001100110111011101110111101110111011101110111011101110111011101110110111001100110011001100110011001011110011001100110011001100110011001100110011001100110011001100110011001101110111011100110111101110111011101110111011101110111011101111111011101101110010111011101110111011101111001100110010111011101010101010101010101010101010101010101110111100110011001101110111101101110010111011101110111011101110111011101111001100110011011101110111011100101110111011101110111011101110111011101110111011101110111011101110111100110011011110111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100101110111011101110101010100110011000100001110111011001100110011101111001110011011100101110111010100101100100001100110011001100100010001000100010001000100011001100110011001100110011001100110011010001000101010101000100010001010101010101100110011110011001100110000110010101000100010001000100010001000100010101100110011110001001101010111100110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011000100010001000011101110111011001100110010101010011001000100001000100010001000100010001000100010001000100010001000100010001000100010010010101100110011001000011000100010001000100010001000100010001001000100010001100110100010101010101010101010101010101010100010001000100,
	2400'b011110001000100110001000100110010111011010000111010101000011001000010001000100010001000100010001001000100010001100110010001100110011001100100010001000100010001000100010001000100011010001000100010001000110100110011001101010101010101010101001100001110111011010000111010101000011001100110011001100110011001100110011010001101001101010111001101010101000011101111000100010011011110011001100110011001011100010000111011101100101010101010110100010111100110111101110111011101110111011101110111011011101110111011100110011001100110011001101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101010000111011101111001100110011000011001100110010101010100010001000100010001010111011110000111011001100110011001110110011110101011110011001100110011001100110111011101110111011110111011101110111011101101110111001100110011001100110011001100101110111100101111001011110010111100110011001100110011001100110011011101110111011101110111101110111011101110111011101110111011101110110111001011101110111011101110101011101010111011101110111010101010101010101010101010101010101010101111001100110111011101110111011101110010111011101110101010101010111011101110111100110011001100110111001100101110111011101110111011101110111011101110111011101110111011101111001100110011011110111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001011110011001011101010101001100010001000011101100101011001110111100110111100101110111011101010000110010000110011001100100010001000100010001000100010001100110100010001000100001100110100010001000100010001000100010001000101011001010111100110011001100001010100010001000100010001000100010001010101011001111000100110011010101010111100110011011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011000100010001001100010001000011101110111011001110110011001010011001000100010001000010001000100010001000100010001000100010001000100010001000100100100011001100110010000100001000100010001000100010001000100010001001000100011001101000101011001100110010101100110011001010101010101010101,
	2400'b011110001000100110011000100110010110011110000110010000110010000100010001000100010001000100010010001000100010001100110011001100110011010000110010001000100010001000100010001000100010001000110011001101001000100110101001101010101010101010101001100001110111011110000111011001000100010001000011001000110011001100110011001101000110100110111010100110111001100001110111100010001001101111001100110111011100101010011000100001110110011001010110011110101101110111101110111011101110111011101110111011011101110111011101110011001100110011001100110011011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111010100101110111100010011001100110101000011101100110010101000100010001000100010001000101100010011000011101100110011101110111011110001011110010111100110011001100110011001100110111011101111011101110111011011101110011001100110011001100110010111011101110111011101110111011101110111011110011001100110011001100110011011101110111011101110111101110111011101110110111101110111011101101110010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101011101111001101110111011101110011001100101110111011101010101010101010101011101110111011101111001100110011001011101110111011101010101011101010101011101110111011101110111011101111001100110011011110111011111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001011110010111011101010011001100110011000100001110110011001100110011010011011101111001011101010011000010100110011001100110010001000100010001000100010001000110011010001010101010000110011001101000100010001000100010001010110010101011000100010000111010101000100001101000100010001000100010101100111100010011001100110101011101110111011110011011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101001100110001000100110011001100110001000100001110110011001010101010101010011001000100010001000100010000100010001000100010001000100010001000100010001000100110101011101100101001100100001000100010001000100010001000100010010001000110100010001010111011101100110011001100110011001100110011001100101,
	2400'b011110001000100010011001100110000110011101110110001100100001000100010001000100010001000100100010001000100010001100110011010000110011001100110010001000100010001000100010001000110011001100110010001101011001100110101010101010101010101010101010100110000111100010010111010101000101010101100100001100110010001100110011001101000100011010101011101010111011100110001000100010001001101011001101110111011100101110101010100110000110011001100101011110011100110111011110111011101110111011101101110111011101110111011100110011001100110011001100110011001101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110010111001100001111000100110011001101010011000011101100101010101010100010001000100010001000101011010011010100110000111011110000111011101111010101110111100110011001100110011001100110011001101110111011110111011011100110011001100110011001011101110111011101110111011101110111011101110111011110011001100110011001100110011011101110111011101111011101110111011101110111011101101110111011100101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101011101111001101110111011100110010111011101110111010101010101010101010101010101010101010101010111011101110111011101110101010101010101010101010101010101010101010101110111011101111001100110111011110111011111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001011110010111010100110011010101010011000100010000111011101100101010101101001101111001011101010101001011101010011001000100010001000100010001100110011001100110011010001010101010100110011001101000100010001000100010001010101011001110111011101100101001100110011001100110011010001000100010101100111100010001001101010101010101110111011110011001101110111011101110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010100110011001100110011001100110001000100010001000011101110111011001100110010100110011001100110011001000100010001000010001001000010001000100010001000100010001001001010110011001010011001000100010001000010001000100010001000100100010001101000101010101010101011101110101010101100110011001100110011001100110,
	2400'b100010001000100110011001100101110110100001110100001000010001000100010001000100010001000100100010001000100010001000110100010001010100010001000011001000100010001000100010001000100011001100110011010001111001100110101010101010101010101010101010100110001000100110010111010101000101011001100110001100110010001100110011001100110011010001101010101110101011101110011000100010001001100110111101110111011101101110111011101010010111011001100101011010001011110011011101111011101110110111011101110111011101110111001100110011001100110011001100110011001100110011001101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110010101000100110101010100110011010100110001000011101100101010101010101010001000100010001000100010101111001101010101010100010001000011101111001101110111100110011001100110011001100110011001100110011011101110111001100110011001100110011001100101110111011101110111011101110111011101110111011110011001100110011001100110011011101110111011101111011101110111011101110111011011100110010111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101111001100110011001100101110111011101110101010101010101010101010101010101010101010101010101011101110111010101010101010101010101010101010101010101010101010101110111011101110111100110011011101111011101111111011111111111111111111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100101110101010101110111010100110011010100110011001100010000111011001010101100010101011100110011010100101110100001100100011001100110011001101000100010001000100010001000100010000110011001101000100010001000100010001010101011001100111011101010011001100110011001100110100010001010110011001110111100010001000100110011010101010101011101111001100110111011100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101001100110011001100110011000100010000111011110000111011101110110011001100110010000110100010101000100001100110010001000100011001100110010000100010001000100010001001001000110010101000011001000100010001000010001000100010010001000100100010101110101010000110011010001010101010101010101010101010101011001100110,
	2400'b100010001000100110011001100101100110011101000010001000010001000100010001000100010001001000100010001000100010001000110100010101010101010001000011001000100010001000100010001000100010001000110011010110001001100110101010101010101010101010101010100110001001100110010111010101010110011101100110010000110011001100110011001100110011001101000110101110111010101110101001100010001000100110101100110111011101110010111100101110101000011101110110011010001010110011011101111011101110110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001101110111011101110011001100110011001100110011001100110011001100110011001100110111011100110010111010101111001011100110011001100001110110011001010101010101010100010001000100010001000100010001010110100110111011101010011001100001111000101110111011110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001101110111011110111011101110110111011101110011001011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111100110010111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011110011001101111011101110111111111111111111111111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100101010111100110010101001101010111010101010101010101010011000011101100100010101111010101001110111011101110101001100100011001101000100010001000100010001000100010001000100010000110011001100110011010001000100010001010101011001100110010100110011001100110011001100110100010101100110011101111000100010001000100110001001101010101011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101001100110011001100110011000100010001000011101110111011001100110011001100110010101000101010101010101010101000011010001000101010101000011000100010010001100100001000101000011010001000010001000100010001000010001000100100010001100110100010001000100001100110010001100110011001100110011010001000100010001000100,
	2400'b100010001001100110011001100001100111011000110010000100010001000100010001000100010001001000100010001000110010001100110011010001010101010001000011001000100010001000100010001000100011001000110100011110011001100110011010101010101010101010101001100010011001100110000111011001100111011101110111010000110011001100110011001100110011001101000100011110111011101110111010100110011001100110011011110111011101110011001100110010101001100010000111011001111010110011011101110111101110110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111001100110011001100110011001100110011001100110011001100110111011101110011001100110011001010100110000111011101100101010101010101010101000100010000110011010001000100010001010101011110011011101110101010100110001000101010111011110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001101110111101110111011101101110111001100101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101111001100110111101110111111111111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011001100101110101011101110101011101110111010100110011000100001110110010101010111100110000101010101110110010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010101000101011001100100001100110011001100110011010001000100010001010101010101100111011110001000100110011010101010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101111001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010011001100110001000100001110111011101110110010101010110011001100101010101010100010001000101010001000011001101000100010001000011001000100010001100110001000100110011010000110010001000100010000100010010001000110011001100110010001000100011001100110011001100110011001100110011001100110011001100110011,
	2400'b100010001001100110001000011101010110010000100010000100010001000100010001000100010010001000100010001000110011001100110011010001010110010001000011001000100010001000100010001000100011001100110110100010011001100110011001100110011001100110011001100010011001100010000111011101110111011110000111010001000011001100110011001100110011001101000100010110001011101110111010100110011001100110101011110011011101110011011101110010111010100110011000011001101001101111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111001100110011001100110011001100110011011100110011001100110111001100110011001100110010111001100001110111011001010110011001010100010001000100010001000100001101000100010101010101010101111001101110111011101110101000101010111011110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001101110111101110111011011101110011001100101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101111001100110111101110111011101110111111101111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011100101111001100110010111011101110111010100110001000011101110111010101000100010101110110010001000100001100110010001000100010001100110011001100100010001000100010001100110011001100110011001100110100010001000101011001010011001100110011001100110011010001000100010001010101010101100110011110001001100110101011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010011001100010000111100001110111011101110110011001100110011001100110010101010101010001000011001100100010001000010001001000100010001000010010001100110001000100100100001100100010001000100001000100010010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011,
	2400'b100010001001100110010111010101100100001000100001000100010001000100010010000100010010001000100010001000110011001100110011010001010101010000110100001000010001000100100010001000100010001101001000100110011001100110011001100110011001100110011001100110011000100010001000011101111000100010000111010101000011001100110011001100110011001100110100010001101010101110111011100110011010100110101011110011011101110011001101110011001100101010011001011101101000101011001101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011001100110011001011101111001100110010101000011001100110011001100111011101010100010001000100010001000100010001000100010101010101010101100111101010111011110010111010101110111011110010111100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001101110111101110110111001100110010111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101111001100110111011110111011101110111111101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110011001010101010101001100010000111011101100110010101000100010001010111011001000011001100100010001000100010001000100011001000100010001000100010001000110011001100110011001100110100010001010110010100110011001100110011001100110011010001000100010001010101011001100110011101111000100110101011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011000011101110111100010000111011101110111011101110110011001100110011001010101010101010100001100110010000100010001000100010001000100010001000100100001000100100011001000100001000100010001000100100010001000100010001000110011001100110011001100110011001101000100010001000100010001000011001101000100,
	2400'b100110001000100001110110010001000011001000100010000100010001000100010010000100100010001100100010001000110011001100110011010001010101010100110100001000100010001000100010001000100010001101011001100110011001100010011001100110011001100110011001100110001000100010001000100010001000100010000111011001010100001100110011001100110011001100110100010001000111101010101010101110101001101010101011110011011101110111001101110111011100101110101010100101100111100111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110011001100110010111100110011001100100110000111011001100110011110001001011001000100010001010101010001000100010001000100010101010101010101010110011110101011110011001011101110111011101111001011110011001100101111001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001101110111101101110011001011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101111001100110011001101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001101110110111011101110101001100110000111011101100110010101010100010001000101011001010011001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011010001010101010000110011001100110011001100110100010001000100010101010101010101100110011001110111100010011010101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010011001100010001000100001110111011101110111011101110110011101110110011001100101010101000100001100110010000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100100010001000100010001000100011001100110011001100110011001100110100010001000100010001000100010001000100,
	2400'b100001110110011001100101001100100010001000100010000100010001000100100010000100100011001100100010001000110011001100110011010001010110010101000100001100100010001000100010001000100011001101101001100110001000100010001001100110011001100110011001100010001000100010001000100010001000100010000111011001010100001100110011001100110011001100110011010001000101011110101010101110111010101010101011101111001101110111011100110111011101110010111100101001110110100010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111001100110011001100110011001001100010000111011001110111100010101000010101000100010101010100010001000100010001000100010101100101010101010101011010001011110011001100110010111011101110111100110011001011110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001011101111001100110111011101101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101111001100110011001100110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011011101110111001100110010101010100110000111011101110110011001100101010101000100010101010100001100100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010101010100001100110011001100110011001100110011001100110100010001010101011001100110011101111000100110101011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110001000100010000111011001100101010101010101010101000100001100110010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001100110011001100110011001100110100010001000100010001000101,
	2400'b011001010110011001100100001000100010001000100001000100010001000100100001000100100011001100100010001101000100001100110011010001010110011001010101001000010010001000110010001000100010001101111001100010001000100010001001100110011001100110011001100010001000100010001000100010001000100010000111011101100100001100110011001100110011001100110011001100110100010101111001101010101010101010101010101111001100110111011100110111011101110010111100101110000110100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011100110011001100110010110111011101110111011101111000101010100110010101000101010101010101010001000100010001000100010001100110011001100101011001111001101111001100110010111011101110111011101110111100101110111100110010111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110010111011101110111100110011001100101110111011101110101010101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111100110010111100110011001101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110011001101110111001100110010101001100110011001100001110111011001100101010101000100010101000100010000110010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010101000011001100110011001100110011001100110011001100110100010101010110011001110111011110001001101010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101001100101110110011001010100010001000011001100110011001100110010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011001100110011001100110011001100100011001100110011001100110011010001000100010001000100010101010101,
	2400'b010101010101011001010011001000100010001000010001000100010001001000100001001000100011001100110010001101000100001100110011001101010110011001010100001000010001001000100011001100100010001101111000100010001000100010001000100010001001100010011001100010001000100010001000100010001000100010000111011101110101010001000011001100110011001100110011001100110100010001100111100110101010101010101010101111001100110111011100110111011101110111001100110010100111011110011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111001100110011001100110011011101110111011101110011011101110011001100110010010110011001110111100110011010101110010101010101010101010101010101010001000100010001000100010001100111011001100110011001101000101010111011101110111011101110111011110010111011101110111011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011110010111100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111001101110111011101110111011101110010111100110011001011101110101000100010011001100110000110011001010101010101010100001100110011001100110011001000100010001000100010001000110011001000100010001100110011001100110010001100110100010000110011001100110011001100110010001000110011010001010110011001100111011101111000100010011001101010101011101111001100110111011101110111011100110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111010101110111011101110101001100001100101010000110011001100110011001100110010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001100110011001100110011001100110011001100110100010001000100010001000100010001010101,
	2400'b010101010110010100110010001000100010000100010001001000100010001000100001001000110100001100110010001101000100001100110100001101010110011001010101001000100001000100100010001100110011010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001110101010001000011001100110011001100110011001100110011010001010110100010011010101010101010101010111011110011011101110111011101110111001100110110111000011110101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110011001100110011001100110111011101110111011101110011001100101001110110011001111000101010101011101101110101010101010101010101010101010101000100010001000100010001100111011101110111011101100111100110111011101110111011101110111011110011001100110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100101110111010101010101011101110111100110111011100101111001100101011001011101010011000100110101010100110000111011001100101010101000100001100110011001100110011001100100010001000100010001000110011001000100010001100110011001100110011001101000100001100110011001100110011001000100011001101000101011001110111011101110111011110001000100110011010101010101011101111001100110011001101110011001100110011001101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110101010101110111010100101110101010000110011001100110011001100110011001100100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000110011001100110011001101000100010001000100010001000100010101010101,
	2400'b011001100101010000100010001000100010000100010001001000100010001000100010001000110100001100110011001101010101010000110100001101000110011001100100001000100010001000100010001000110011010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110010001010100001100110011001100110011001100110011001101000101011110011010101010101010101010111011110011001100110111011101110111011100110111001001100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011100110011001100110111011101110111011101110011001011011101100110011010001010101111001011100101100101010101010101010101010110010101000101010101000100010001010111100010000111100110000110100010101011101110111011101110111011110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101111001100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110011001011100110011000100010001000100010001001100110011000101010111010101010011001011001010110011001110111011110001000011101100101010101000100010000110011001000100010001000110010001000100010001000110011001000100010001000110011001100110011001100110011001100110010001100110010001000110011010001010110011001110111011101111000100010011001100110011010101110111011101110111011101111001100101110111100110011011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111010101110111010101010000110010000110011001100110011001101000011001100110010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011001101000100010001000100010001000100010001010101010101010101,
	2400'b011001010101001100100010001000100010001000010010001000100010001000100010001001000100010001000011001101010101010001000101010001000110011001100100001000010010001000100010001000100011010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100001110101010101100100001100110011001100110011001100110011001101000100011010001010101010101010101010101010101111001100110011001101110111011100110111001010101010101011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110011001101110111011101110111011101110010111000011001100110011110011011101111001011100001100101011001100101010101010110010101000101010101000100010001010110100010011000101010100111011110011011101110111011101110111011110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101111001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011100101110111011101010011000100001110111011101110111011001100110011001100110011101100110010101010100001100110010001101000101011101110111011001000100010001000100001100100010001000100010001000100010001000110011001000100010001000100010001100110011001100110011001100110011001000100010001101000100010101100110011001100111011110001001100110011001100110101011101010011000100010101011101111001100110011011101110111011101110111011101110111011100110011001100110011001100110011001100110011001101110111011100110011001100110011001100101110111011101110111011101110111011101110111011101110111010101110101000011001000011001100110011001100110100010000110011001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100110011010001000100010001000101010101010101010101010101,
	2400'b011001010100001000100010001000100010001000010010001000100010001000100010001001000101010001000100010001010101010101000101010101000101011001010011001000010001001000100010001000110011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100001110101011001110101001100110011001100110011001101000100001100110100010101111001101010101010101010101010101011001100110011001101110111011100110111011011101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111001101110111011101110111011101110010010111011101100110011110101100110011001010011101100110011001110110010101010110010101000101011001010100010001010110100010011000100110111001011110001010101110111011101110111011110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101111001100110011001100110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101111011101101110111001100110010111011101110011001100110011000100010000111011001100111011001110110011001100101010001000100010000110011001000100010001101000110011001010100001101000100010000110011001000100010001000100010001000100010001000100010001000100010001101000011001000100011001100110010001000110011010001000101010101010110011110001001100110011001100110011001100110011000011101111000100110101010101110111100110011001100110011001100110011001100110111001100110011001100110011001100110011001100110111011101110111011101110011001100110011001100101110111011101110111011101110111011101110111011101110111010100001100100001100110011001100110100010001000011001100110011001000100010001000100010001000100010001000110100001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000110100010001010101010101010101010101010101010101010101,
	2400'b010101000010001000100010001000100010000100010010001000100010001000100010001101000101010001000100010001010110010101000101010101000101011001010011001000100001000100010010001000110101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100001110110011101110101001100110011001100110011001100110100010000110011010001011000101010111011101010101010101010111100110011001100110011001100110011011011101010101010101111001100101111001100110011001100110011001100110011001011110010111011101110111011101110111100110011001100110011001100110011001100110111011101110111011101110111011100110111011100101001110110011101110111100010111100110010111000011001100110011101110110010101010101010101010110011101010100010001010110100010011000100010111011100010001001101010111011101110111011110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101111001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011100101110111100110010111011101010111010101010101001100010000111011110000111100010000111011101110101010101010110010101000100001100110010001000100011010001010100010001000100010001000100001100100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001100110011010001000101011101111000100110101001100110000111011101100110011001010101010101100111011110001000100110011010101010101011101110111011110011001100110011001100110011001100110011001100110011001101110111011101110111011101110011001100110011001100101110111011101110111011101110111011101110111011101110100111010000110011001100110011010001000100001100110011001000100010001000100010001000100010001100100010001000110100010000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010101010110011001010101010101010101010101010110,
	2400'b010100110010001000100010001000100010001000100010001000100010001000100011001101000101010101000100010001010110011001000101010101010100011001010011001000100010001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100001100111100010000101001100110011001100110011001100110100010001000011010001010110100110101011101010101010101010111100110011001100110011001100110011001011101110101001101110111011101111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011110011001100110011001100110111011101110111011101110111011101110111011011100001110111011110001000100110111100110010101000011001100111100010000110010101010101010101010111100101100101010101010110100010101001100010111100101010001000100110111011101110111011101111001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101111001100110011001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011100110011001100110010111011101111001011101110111001100110001000100010001000101010011001101010010111011110000111010101010110010101010100001100100010001000110100010101010100010101010101010000110010001000100010001000100010001000100010001000100010001000110011001000110010001000100011001100110100010101101000100110011001100001110101010101000011001100110011001100110100010001000100010101010110011001110111011110001000100110101010101110111011110011001100110011001100110011001100110011001101110111011101110111011101110111011100110011001100101110111011101110111011101110111011101110111011100101100100001100110100010000110011001100110011001100110011001100110011001100100011001100110011001100110010001100100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001101000110011001100110011001100110011001100110,
	2400'b001100100010001000100010001000100010001000100010001000100010001000100100001101010110010101000101010001010110011001010101010101010100010101010011001000100010001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000011101101000100010000101010001000011001100110011001100110011010001000011001101000101100010101011101110101010101010101011110011001100110011001100110011001011101110101001101110111011101110111011110010111011101110111100110010111011101110111011101110111011101110111011101110111011110011001100110011001100110011011101110111011100110011011101110010111000011101110111100010001001101010111100101110011000011001100111100010010111010101010101010101011000100101110101010101010110100010101001100010101100110010011000100010101011101110111011101110111011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001101010101010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101111001100110011001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111001100110011001100110010111100110011001100110010101001100110011001100110011010101110101010101010001000011101110110010101100110011001100110010100110010001000100010010001010110011001010110010101010100001100100010001000100010001000100010001000100010001000100010001000110010001000110011010001010111100010001001100101110101010000110011001000100010001000100010001100110011001100110011010001000101010101100110011101110111100010011010101010111011110011001100110011001100110011001100110111011101110111011101110111011101110111011100110011001100101110111011101110111011101110111011101110111010011001000011010001000100001100110011001100110011001100110011001100110011001100110100010001000100010000110011001100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100100010101100111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001100100010001100110100010001010110010101010101010001010110011101100100010101100101010101010010001000100010001000100011001101011000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100110001001100110001000011001111000100010000101010101000011001100110011001100110011010001010100001101000100011010011010101110111011101010101011110011001100110011001100110011001011101110101001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001101110111011101110011001100110010010111100010001000100110011010101110111100101010101000011001111000100110101000011001010101010101101001101010000110011001100111100010111010100010001011110010111000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001101010011010101010101001100110101010101010101010101010101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011110011001100110011001100110011001101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011100110011001100110011001100110011011100110011001100110011001100101110101010101010101010101010101100110010101001100001111000011101110110011001110110011001100110011001010100001100100010001000110101011101110111011001100110010100110010001101000100001100100010001000100010001000100010001100110010001000110100010101111000100001110101010000110011001000100010001000100010001000100011001100110011001100110011001100110100010001010110011001111000100010011010101010111011110011001100110011001100110011011101110111011101110111011101110111011101110111011100110011001100101110111011101110111011101110111011101010100111010000110100010000110011001100110011001100110011001100110011001101000100010001010101010101100101010101000100010000110011001000100010001000100010000100010001000100010010001000100010001000100010000100010001000100010010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001101010110011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001100100011010000110100010001010110010101010101010101010110011101100101011001100110010101000010001000100010001000110011010001101000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000100010000111011110001000100001110101011001010100001100110011001100110100010001000100001100110100010110001010101110111010101010101011110011001100110011001100110011001011101110101001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001101110111011101110011001100101010001000100110001010101110011011110010111011101010111000011110001001101010111000011001010101010101111011101110010111011101101000100110101011100010001010110011001010100010011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001101010101001100110101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110011001100110011001100110011011100110011001100110011001011101010111011101110101010101010101011101110101001100110101001100010011001100001110111011101100101010101100110010101000011001100100010010001111000011110001000100001100011001001100111010000110011001000100010001000100010001100100011010001000101011001100110010100110011001000100010001000100010001000100010001000100010001000110011001100110011001100110011010001000101011001111000100110101010101110111100110011001100110011011101110111011101110111011101110111011101110111011101110111011100110011001100110010111011101110111011101110111011101001100100001101000100001100110011001100110011001100110011001100110100010001000101010101100110011001110110010001000100010001000100010001000100010000110011001000010001001000100010001000100010001000100001000100010001000100010010001100100001000100010001000100010001000100010001000100010001000100010001000100010001001000100100011010001000100010001000,
	2400'b001000100010001000100010001000100010001000100011001100100011010001000100001101000110011001010101010101010110011101110110011001100110011001000010001000100010001000110100011010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110001000100010000111100010001000100001110101011001010101001100110011001101000100010001000101010000110100010101101001101010111010101010101011101111001100110011001100110011001011101110111001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001010100010011010101110101011101110101010101110111011101110111001011110001001101110111001011001100110011010011011101110011000011101101000101010101011100110001001101111001011100110011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110101001100110101001100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101111001100110011001100110011001100110011001100110111101110111011101110111011101110111011101110111011101110111011101110111011101101110111011100110011001100110011001100110011001100110011001100110011001100110010111010101111001011101110101010101010101011101010011001100010000111011101110111011101100101011001010110011001100110011001100110010100110010001000110110100010001001101010010110001001011000010101100110010001000010001000100010001000100011010001010101010101000011001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000100010101010111100010011010101010111011110011001100110011001101110111011101110111011101110111011101110111011101110011001100110011001100110010111011101110111011101110111010011101000100010001000100001100110011001100110011001100110011010001000100010101010110011101110111011101110111010100110011001100110011001101000100010000110010000100010001000100100010001000100010001000010001000100010001000100010011010000110010001000110010001000100010000100010001000100010001000100010001000100010001000100010010001101010110100010001001,
	2400'b001000100010001000100010001000100010001000100011001100110100010101000100001101000110011001100101010101010110011101110110011001100110011001000010001000100011001100110101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000100001111000100010001000100001100110011001100110010000110011001101000100010001000100010101000100010001010111101010111011101010101011101110111011110011001100110011001011101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110010101001101010111011101110111100101110011010101110111011101110111001011110011010101110111010011101100111100110111100110010101000100001111000101010101011101010001001101010111100101010011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101001101010011001100110011010100110101010100110011001100110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101111011101110011001100110011001100110011001101110111101110111011101110111011101110111011101110111011101110111011101110111011101101110111001100110011001100110011001100110011001100110011001100110011001100110010101010110011001011101110111011101010011000011101100101010101010100010001010100010001000100010001010101010101010101010101100110011101100101010000110010010101111001101010011000001100110111010101111000011101110011001000100010001000100011010000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110100010001000100010001000101011010001001101010111011101111001100110011011101110111011101110111011101110111011101110111011101110011001100110011001100101110111011101110111011101110100111010001000100010000110011001100110011001100110011001100110100010001010110010101100111011101110111011101110111011001000011001100100010001001000100001100100001000100010001000100010001000100010001000100010001000100010001000100010010010000110011001101000011001100110011001000010001000100010001000100010001000100010001000100010001000100100011010110001001,
	2400'b001000100010001000100010001000100010001000110011001100110100010101000101010001000110011001100101010101100110011101110111011001110111011001010010001000100011010001000101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100111011101110110010000110011001101000100010101010100010001010100010001010110100010101011101010011010101110111011101111001100110011001011101110111010101010111011101110111011101110111011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101110111100110011001011101110001010101110111011101110111010011110011010101110111010011101101000101111001100110010111001100001111000101010111100101110011010101010111100101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101010100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011110011011110110111011100110011001100110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111001100110011001100110011001100110011001100110011001100110011001100110010111100110011001011101010011000011001010101010101010101010101010101010101010101010101010101010101100110011001100110010101010101010101010111011101100100001000110111100110101001010100100101010001100111011101000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100100011001100110011001100110011001100110100010001000101010101010101010101010111100110101010101111001100110111011101110111011101110111011101110111011101110111011100110011001100110011001100101110111011101110111011101001110100010001000100001100110011001100110011001100110011001101000101010101010111011101100111011101110111011001100110010101010011001100100010001001000100001000010001000100010001000100010001000100010001000100010001000100010001000100010010010000110100010001000100010000110010001000100010000100010001000100010001000100010001000100010001000100010010001101011000,
	2400'b001000100010001000100010001000100010001100110011001100110101010101000101010001000110011001110110010101100110011101110111011001110111011001010010001000100011010101010110100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111010000110011001100110100010001010100010001010101010001010101011010011011101010101010101110111011101110111100101110111011101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001011101010001010101110101011101110101010100010011010101110111010011101111010110011011101110010111001100010001001101010111011101110101010101010111100101110111011101110111011101110111011101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001101110111001100101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011010100110011010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111100110111101110111011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101001011101100110011001010101010101010101011001010101010101010110011101110111011110001000100010001000011101110111011001010101010101100110010000100011011010011000010100100011001101000110001100100010001000100010001000100010001000100010001000100011001100100010001000110011001100110010001100110011010001000100010001000100001100110011001100110011010001000100010101010101010101010101011010001010101111001100110111011101110111011101110111011101110111011100110111001100110011001100110010111011101110111011101110111010011101000100010001000100001100110011001100110100001101000100010001010111100001111000011101111000100010001000100001110101010000110011001000100010001000110011001000010001000100010001000100010001000100010001000100010001000100010001000100010010010001000100010101010100001100100001001000110010000100010001000100010001000100010001000100010001000100010001001000100100,
	2400'b001000100010001000100010001000100010010000110011001100110101010001000101010001000101011001110110011001100111011101110111011001110111011101100011001000100011010001010111100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011110000111010100110011001100110100010001010101001101000101010101010101010101111010101010011010101110111011101110111011101110111011101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110010111011100110001010101010101010101010101010100110011010101110111001011110011100110011011100110010111001100010001010101110111011101110111011101010111011101110111011101110111011101110111010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001101110111011110111011101101110110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101111001101111011101110111011101110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001011100101110111011001100110011001100110011001100110011101100110010101100111100110011010101010101010101010101001100110101010100110010111011001010101010101000010001001000110010100100010001000110011001000100010001000100010001000100010001000100010001000100011001100110011001101000100010000110011001101000100010101100110011001010110010101010100010001000100010001000100010001010101011001010101010101101001101111001101110111011101110111011101110111011101110111011100110011001100110011001100110010111011101110111011101110100111010001000100010001000011001100110011001100110101010001000101010001011000100110011001100010001000100110001001100010000111010100110011001000100010001100110010001000010001000100010001000100010001000100010001000100010001000100010001000100010011010101010101010101000011001000010010001000110010001000100001000100010001000100010001000100010001000100010001000100010010,
	2400'b001000100010001000100010001000100011010000110011001101000101010001000110010101000101011101110111011001100111011101110111011101110111011101100100001000100010010001011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010000111010101000011001100110100010001010101010000110100010101010101010101101000101010101010101110111011101110111011101110111011101110111010101010111011101110111011101110111011101110111010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011010101010101010101010101010100110011010101110111001100010101100110011001100110010101001100110011010101110111011101110111011101110111011101110111011101110111011101110101010101010101010101110111011101110111011101110111011101110111011101110111100110011001100110010111011101110111011101110111011101110111011101110111011101111001101111011101110111011011101110111001010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101001100110101001100110011001100110011001100110011001100110011001100110011001101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010111011110011001011110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110011001100110011001100110011001100110011001100110011001100101110101000011101110111011001110111011001111000011101111000100110000111011110001001101010111100110011001011101010011001101010101010101010011001101010011000011101010011001000100011010000100010001000100010001101110101001000100010001000100010001000100010001000100010001100110011001100110100010101000011001101000101010101100111011101110111011101100110011001010110010101000100001101000100010101100110010101010110100111001100110111011101110111011101110111011101110011001100110011001100110011001100110011001011101110111011101101110100010001000100010000110011001100110011001101000101010101010101010101010110100110101001100110011001100110001000011101100110010101000011001000100010010000110010001000010001000100010001000100010001000100010001000100010001000100010001000100010011010101010101010000110010001000100010001100100011001100100001000100010001000100010001000100010001000100010001000100010001,
	2400'b001000100010001000100010001000110100010000110011001101000101010001000110011001000101011001110111011101100111011101110111011101110111011101110101001100110011010001101001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010000111011001010100001100110011010001000101010000110100010101010110011001010111100110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100010011010101010101010101010101010101010011010101110111001100010101011110011001100101110101001100110101011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101011101110111011101110111011101110111100110011001100110011001100110011001100101110111011101110111011101110111011101110111011110011011101111011101110111011101110110111001010101010101010101010101010101010101010101010101001100110011001101010101010101010101010101010101001100110011001100110011001101010101001100110011001100110011001100110011001100110011001100110011001101010011001101010101010101010101010101010101010101010101010101010101011110011001100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110011001100110011001100110011001100110011001100110011001011100110000111011101111000011101111000011110001001100110011010101010011001100110011011110011001100110010111010101010011001100010000111011101100110011001100111100010000110001100100010001000100010001000100011100010010101001000100010001000100010001000100010001000100010001000100011001100110100010101010100001101000101011001110111011101110111100001110111100010000111011101100101010001000100010001010101011001010101011110101100110111011101110111011101110111011101110011001100110011001100110011001100110011001100101110111011100001010100010001000100001100110011001000110011001101000101010101010101011001100110011110101010101010101001100110000111011101100101010100110011001100100011001100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010011010101010100001100100011001100110011001100110011001100100010000100010001000100010001000100010001000100010001000100010001,
	2400'b001100100010001000100010001000110101010001000011001101000101010001010110011101010100011001110111011101110111011101110111011101110111011101110101001100110011010101111001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001111000100010001000100010000111011001100100001100110011010001000110010101000100010001010110011001100110100010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100010011010101010101001100110011001101010101010101010101000100110101011101110111100110010111010101010101011101110111011101110111011101010111011101110111011101110111011101110101010101010101010101010101010101010101010101010101011101111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111100110111011101110111011101110111011101110111001011101010101010101010101010101010101010101010011010100110011001100110101010101010101010101010101010100110101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010111100110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110011001100110011001100101110101001100010001000100010001000100010011001100110011010101010111011101110101011101110111100110011001011101010000111011001100101010101000100010000110011001100110011010001100111011000110001001000100010001000100101100110000100001000100010001000100010001000100010001000100010001000100010001000110011010001010101010001000101011110001001100110001000100110000111100110011000100110010111010101101000011101100101011001110111011110001010110011011101110111011101110111011101110111001100110011001100110011001100110011001100101110111001010101000100010001000100001100110011001100110011010001010101010101010110011101111000100010001010101010101001100110000111011001100110010101010011001100110011001100100010001000010001000100010001000100010001000100010001000100010001000100010001000100100100010101010100010001010100010001000100010000110011001100100010001000100010001000010001000100010001000100010001000100010001,
	2400'b001100110011001000100010001001000101001101000011010001010101010001010110011101100100011001110111011101110111011101110111011101110111011101110101001100110011010101111001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010000111011101110101010000110100010001000110010101000100010001010101011101100110011110011010101010101010101010101010101010101010101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100010101010101010101001100110011001100110101010101010101001100110101010101110111100110010111011101110111011101110111011101110111010101010111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111100110111011101110011001011110011001100110011001011101010101010101010101010101010101010101010011001100110011001100110101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101011110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110011001100110011001011100110011001100010001000100110011001101010101010101010101011101110111011101110111011110010111011101010011000011001010101010000110011001100110010001000100010001000100010001000110011010101110100001000100001001000100011010100110010001100110011001000100010001000100010001000100010001000100010001000100011001101000100010001000110100010011001101010101001101010101001100110101010101010101010100010001010101110011000011110011011101010001000101111001101110111011101110111011101110111001100110011001100110011001100110011001100110010010101010001000100010000110011001100110011001100110100010001010101011001100111011110001001100110011001101010101001100110000111011101110111011001010011001100110011001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100100101011001100110011001010101010101010100010001000011010000100011001000100010001000010001000100010001000100010001000100010001,
	2400'b001100110011001000100010001101010101001101000100010001010101010001010110011101110101011001110111011101110111011101110111011101110111011101110100001100110100010110001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110101010001000100010001000110011001000100010001000101011001110110011010011010101010101010101010101010101010101010101010101011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100010101010101010011001100110011001100110011010101010011010101010101010101010111011110011001011101110111011101110101010101110101010101010101010101110111011101110111011101010101010101010101010101010101010101010101010101010101010101111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111101110111001011101010101010101110111011101110101010101010101010101010101010100110101010100110011001100110011001100110101010101010101010101010101010101010101001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110101010101010101010101010101010101010111011110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110011001100110011001100110010111001100110011001100110011001101010101010101110111010101010111011101110111011101010101011101010011001011101010101010001000100001100110011001000100010001000100010001000100010001000100010001001000110001100100010001000100010001000100100011001010101010001000100010001000100010000110011001100100010001000100010001000110011001100110101011010001000100110101010101010101010100110101010101010111011101110111011101110111011100110011011110010111001100010111100110111011100110111001100110011001100110011001100110011011100110111001100101001100100010001000100001100110011001100110011010001000100010101010110011001100111100010011010100110101010100110011001100010001000011101110111011001010011001101000011001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010100011001100110010101010110011001100101010101000100001100110011001100110011001000100010000100010001000100010001000100010001,
	2400'b001100110011001000100010010001100101010001000100010001100101010001100110011101110110010101110111011101110111011101110111011101110111011101110100001100110101011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110101010101000100010001000101011001000100010001010101011001110111011010001001101010011010101010101010101010101010101010101011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111000100010101010101010011001100110011001100110011010100110011010101010101010101010101011101111001011101110111011101010101010101010101010101010101010101010101010101010111011101010101010101010101010101010101010101010101010101010101011101111001100110011001100110011001100110011001100110011001011101110111011101110111010101010111100101110101010101010101010101010101010101010101010101010101010101010011001101010101010100110011001100110011001100110101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110101010101010101010101010101010101010101011110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110011001100110011001100110010101001100110101010101010101010101010111011101110111010101010111011101110101001100010001000011101100110010101010101010001000011001100100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001000100101011010001000011101010101010101000101010101010100010001000011001100100010001000100010001000100011010001000101011001111000100110011001100110101010101010101011101110111011101111001011101110111100110011001011100110001010110011001100110011001100110011001100110011001100110111011100110011001011011101000100010001000011001100110011001100110100010101000101011001100110011101111000100110011010101010101010100110011000100010001000100010001000011001000011001101000011001000100010000100010001000100010001000100010001000100010001000100010001000100010001001000100100011001100110011001100110011001100110010101010100010001000011010001000100001100110010001000010001000100010001000100010001,
	2400'b001101000011001000100011010001100100010001000100010101100101010001100110011101110111010101110111011101110111011101110111011101110111011101100011001101000101011010011000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010001000011101110110010101000100010001000101011001010100010001010110011001110111011001111001100110011001101010101010101010101010101010101011101110111011101010101010101010011001100110011001100110011001100110101010101010101010101010101011101110111011101110111011101110101010101010101010101010111011101110101010101110111011101110101000100110101010100110011001100110011001100110011001100110011001100110011010101010101011101111001100101110111010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101011101111001100110011001100110011001100110011001011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001101010011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101111001101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001101110111011101110111011101110010101010101010111011101110101010101110111011101110101001100110011000100001110110011001100110011001010101010101010101010001000011001000100010001000100010001000100010001000110010001000100010001000100010001000010010001000100010001000100011010101111000011101010100001100110011010001000100010001000100010000110011001000100010001000100010001000110011001101000100010101100111100010011010101010101010101110111011101110111100110011001100110011001100101110011001101011001100110011001100110011001100110011001100110111011100110010110111010001000100010001000011001100110011001101000101011001010101011001100111100010001001100110101010101010101010100110011000100010001000100010011000011101000011010101010011001000100010000100010001000100010001000100010001000100010001000100010001000100010001001000100101011001110111011101110111011001100110011001010101010101000100010001010100010001000011001000100010000100010001000100010001,
	2400'b001100110011001000100011010101100100010001000100010101100101010001100110011101110111011001100111011101110111011101110111011101110111011101100011001101000101011110001000100010001000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011000100010011001100010001000100010000111100001110110011001000100010001010110011001010100010001010101011001110111011101101000100110011001100110011001100110011001101010101010101110111010101010101010100110011001100110011001100110011001100110011001101010101010101010101010101010101011101110101010101010101010101010101010101010101010101010011010101010111011101110101000100110101010100110011001100110011001100110011001100110011001100110011001101010101011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011010101010101010101010101010101010101010101010101010101111001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011100101110111011101110111011101110111011101110111010100110000110011001100110011101100101010101100110010101010101010101010101010000110010001000100010001000100010001000100010001000110011001000100010001000100010001000010001001000100010001000100010001000110011001100100010001000100010001000100010001100110100010001000100001100110010001000100010001000100010001100110011001100110100010101101000100110101010101110111011101110111011110011001100110011001100110010111010101010111100110011001100110011001100110011001100110011011101110010000100010001000100010001000011001100110011010001010101011001100101011001110111100110011001100110101010101010101001100110001000100010001000100010011000011000110011011001000011001100110010000100010001000100010001000100010001000100010001000100010001000100010001000100100100011001110111011101110111011101110110011001100110011001010101011001100101010101000100001000100010001000100001000100010001,
	2400'b010000110010001000100011010101010100010001000100011001100101010101100110011101110111011001100111011101110111011101110111011101110111011101010010010001000101011110001000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100110011000100010001000100010001000100010000111011001010100010101010110011101010100010001010101011001110111011101100111100110011001100110011001100110011001100110101010101010101010101010011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010111010101010011000100110101001100110011001100110011001100110011001100110011001100110011001101010101010101110111011101110111011101010101010100110011001101010101010101010101001101010101010101010101010101010101010101010101010101010101010101010101011110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111010101010101011101110101010101010101010101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010111100110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011100101110111011101110111011101110111011101010011000011001100101010101111000100001110111011101100101010001010101010101010101001100110010001000100011001000100010001000100010001000100011001000100010001000100010001000100001001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000110011001100110011001100110011001000100010001100110011001100110011001101000101011001111000101010101011101110111011101110111011110011001100110011001011101110111010110011001100110011001100110011001100110011011100100101010100010001000100001100110011001101000100010101100110011101110110011110001000100110101010100110101010100110011000100010001000100010001000100010000111010000110011010101000100010000110010000100010001000100010001000100010001000100010001000100010001000100100010001000100011010101100111011101110111011101110110011001100110011001010110011101100110010101010100001100100010001000100001000100010001,
	2400'b010000110011001000110100011001010100010101000100011001110100010101100110011101110111011101100111011101110111011101110111011101110111011101000010010001010101100010001000100010001000100010011001100110011001100110001000100010001000100010001000100010001000100010001001100110011001100110011001100010001001100110001000100010001000100010000111011101010101010101010110011001100100010001010111011101110111011101100111100110011001100110011001100110011001100110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010101010101010011000100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010100110011001100110011010101010101001100110011001100110101010101010101010101010101010101010101010101010101011101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010111100110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101111011011101110111001011101111001011101110111011101010101001100001110110010101010101011110001001100110011001011101000100010101010110010101010100001100100010001000100010001100110011001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000100100011001100110010101000010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001101000101011110011010101110111011101110111011110011001100110011001100110010111010101111001100110011001100110011001100110011001010010101000100010001000100010001000011001101010101010101100111011101110111011110001001101010101010101010011001100110011001100010001001100110011001100110010111010000110011011001100101010000110010001000010001000100010001000100010001000100010010001000100010001000100011001000100011001101010110011101110111011101110111011101100110010101100111011101100110010101010100001100110010001000100010000100010001,
	2400'b010000110011001100110100011001100101010101010101011001100101011001110110011101110111011101110111011101110111011101110111011101110111011000110010010001010110100010001000100010001000100010001001100110011001100110001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100010001000100010001000100010001000011101010101010101100110011001100100010001010111100010000111011101100110100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101000101010101010101010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010111011101110111011101010101010101010111011101110111011101110111011101110111011101110111011101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011110011011110110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011110111011101101110111001100110011001100110010111011100110000111011001100110010101100111100010011001101010010111010101000100010101010110010101000011001100100010001000100011001101000100001100110011001100110011001000100010001000100010001000010010001000100010001000100010001001001001101010101001100001100011001000100010001000100010001000100010001000100010001000100011010001000100001100110011001100110011001100110011001100110011010101101001101010111011101110111011101110111011110011001100110011001011101111001100110011001100110011001100110010110110010001000100010001000100010001000100010001010101011101110111011101110111100010011010101010101010101010101001100110011001100110011001101010101010101010101000010000100101100001110100010001000011001000010001000100010001000100010001000100100010001000100010001000110011001100110011010001010110011001110111011110000111011101100111011101110111011101100101010101010101010000110011001100100010001000100001,
	2400'b010000110011001100110100011001100101011001100101011001110101011001110111011101110111011101110111011101110111011101110111011101110111011000100010001101010110100010001000100010001000100010001001100110011001100110011000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100010001000100010001000100010001000011101100110011001100110011101100100010001000110100010011000011101100110100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010001000101010101010101010010111100110101010100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010100110011010101010101010101010011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101011101110101010101010011001101010101011101110111011101110111011101110111011101110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111101110111011101101110111001100110011001100110010111010100110001000011101110111011001111000100110011010101001110100010001000100010101010101010100110011001100110010001100110011010001000101010001000100001100100010001000100010001000100010001000100010001000100010001000110011001100110110101110111011100101010011001100100011001100100010001000100010001000100010001000100010001000110011001101000011001100110011010001000011001100110011010001010110100110101011101110111011101110111011101111001011101111001100110011001100110011001100110011001100110001110100010001000101010001000100010001000100010101010110011101110111100010001000100110101010101110111011101110111010100110011001100110101010101010101010101010101000010000110110100001100011010000110010000100010001001000100010000100010001000100010010001000100010001100100010001100110011010001100110011101111000100010001000100010001000100001110111011101100101011001010101010001000011001100110011001000100001,
	2400'b001100110011001100110101011001100101011001100110011001100101011001110111011101110111011101110111011101110111011101110111011101110111010100100010001101010111100010001000100010001000100010001001100110011001100110011001100010001000100010001000100010011001100110011000100110011001100110011001100110011001100010001000100010001000100010001000011101100110011001100110011101100100010001000101100010011001100010000111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011000100010101010101010100111100010101010100001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011001100110011001100110101010101010111011101110111011101110111011101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101110111010101010101010101010101010101010101010101010101010101010101011101111001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111101110111011011101110111011101110111011100110010111010100110011001100010001000011110001001101010101010100001000100010001000100010101010101010000110011010000110011001101000100010001010101010101000100001100100010001000100010001000100010001000100010001000100010001000110100010000110011100011001100100101100100001100110011001100110011001000100010001000100010001000100010001000100010001000110011001101000100010001000011001100110011001101000100011010011011101110111011101110111011101110111011101110111100110011001011110011001100110011001100100101010100010001010100010001000100010001000100010101100110100010000111100010011001100110101011101110111010101110111011101010011010101010101010101010101010101010101000001100110111100001000011001100100001000100010001001000100010000100010001000100010001001000100010001000100011001100110011001101000110011101110111100010001000100010001000100010000111011001100111011001100110010101000011010000110011001100100010,
	2400'b001100110011001101000101011001100110011001100110011001100101011001110111011101110111011101110111011101110111011101110111011101110111001100100010001101010111100010001000100010001000100010011001100110011010100110011001100110001000100010001000100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100001110111011101100110011101100100010001000101011110011001100110011000011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001001101010100111011110011001011110001001100110001001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010100110011001100110011001100110011010101010101011101110111011101110111011101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010111011101110111010101010101010101010101010101010101010101010101010101010101011101111001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011100110010111010100110011001100110011000100010011001101010010111010001000100010001000100010101010100001100110100010001000011001101000100010001010110010101000011001000100010001000100010001000100010001000100010001000100010001000110100010001000011010010011100101001100100001101000011010001000011001100100010001100100010001000100010001000100010001000100010001000110100010001000011001100110011010000110100010001111010101110111011101110111011101110111011101110111011101110111011101110111100110011001011011001000101010101010100010001000100010101010101011001100111100010001000100010011001101010111011101110111011101110111011101010101010101010111010101010101010101010100111001100111000011101000011001000010001000100010001001000100001000100010001000100100010001000100010001000100010001100110011010001000101011001110111011110001000100010001000100010000111011001110111011101110110011001000100010001000100001100110010,
	2400'b001100110011001101000101011001100110011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110110001000100010001101101000100010001000100010001000100010011001100110011010101010101001100110001000100010011001100110011001100110011001100010011001100110011001100110011001100110001000100010001000100010001000100010000111011101100111011101100100010001000101011110011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100110010111011110011000011110001000011101111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010011001100110011001100110011001100110011001101010101011101110111011101110111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011101110111011101110111010101010101010101010101010101010101010101010101010101010101011101111001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111001100110011011101110111011100110010111010101010101010101010001000100110011001100101100100001101000100010001000011010001010100001101000100010101010100001101000101010001010110010100110010001000100010001000100010001000100010001000100010001000100010001000100011010001000100001101001001101001110100010101000100010001000011001000110100001100100010001100110011001000100010001000100010001000100010010001000100001100110011010001000100010001010111101010111011101110111011101110111011101110111011101110111011101110111011110010111000010101010101010101010100010001000100010101010110011101110111100010011001100110011010101010111011101110111011101110111011101110101010101110111010101010101010101110100111001101001000010100110011001000010001000100010001000100010001000100010001000100100010001000100010001000100010001000110100010001010110011001110111011110001000100010001000100001110111011101110111011101110110011001010101010001000100010000110011,
	2400'b001100110011001101010101011001100110011101110111011001110110011101110111011101110111011101110111011101110111011101110111011101110101001000100010001101101000100010001000100010001000100110011001100110101010101010101001100110011001100110011001100110001000100010001000100010011001100110011001100110011001100010001000100010001000100010001000100010001000011101110111011101100100010001000100011010011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011110001001100010010111011010000111011110000111011001110111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011001100110011001100110011001100110011001100110011001101010101010101110111011101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011101110111100101110111010101010101010101010101010101010101010101010101010101010111011110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111001100110011001101110011001100110010111011101110111010100001010111100110011000011001000100001101000100010001000011010001010101010001000100010001010110010000110101010001000100001100110011001000100010001000100010001000100010001000100010001000100010001000100010010001010100010000110100100010000110010101010101010101010100010001010101001100100011010000110011001100100010001000100010001000100010001000110100010000110011001101000100010001000101011110101010101010111010101010111011101110111011101110111011101110111011101110100101010101010101010101010100010001010101011001100111011101111000100110011001100110101010101110111011101110111011101110111011101110111011101110111011101110101010101110100110001101010111010000110010001000010001000100010001000100100001000100010001001000100010001000100010001000100010001000110011010101010110011101110111100010001000100010001000100010000111011101110111011001100110011001100110010001010100010000110011,
	2400'b010001000100010001010101011001100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110011001000100010001101101000100010001000100010001001100110011001101010101010101010101010100110011001100110011000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010001000100010001000011001111000011101100101010001000101011010001001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000011101111000100010000110010101110110011101110110011001100111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011101111001100101110111011101010101011101110111010101010101010101010101010101110111011110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111001100110011001100110011001100110010111011101110101001010101000101011001110110010001000100001100110100010001000100010001000101010101010101010101010110011001000100010000110010001100110011001000100010001000100010001000100010001000100010001000100010001000100010001001000101010101000011010001110111011101110110011001010101011001100101010001000101010001000011001100110010001000100010001000100010001000100011010001010100001101000100010001000100010001111010101010101010101010111011101110101011101110111011101110111011101101110101010101010101010101010101010001010110011001110111100010001001100110011010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110100101001101010110010000110010000100010001000100100001001000100001000100010001000100100010001000100010001000100011001100110011010001010110011101111000100010001000100010001000100001110111011101100110011001100111011101100110010101100101010000110011,
	2400'b010001000100010001010110011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101100010001000100010001101111000100010001000100010011001100110101010101010101010101010101010101010101001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000011101100101010001000101011010001001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101110111100010000110010001010110011101100110011001100111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011101110111011101110111011101010111100110010111011101110101010101010111011101110111100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111001100110011001100110011001100110010111011101010010110010000110011010001010100010001000100001101000100010001000101010101010110011001100101011001100110011001000011001000100010001100110011001000100010001000100010001000100010001000100010001000100010001000100010000100100100010101010100001101001000100010000111011101100111011101100101010101100101010101000100010001000011001100100010001000100010001000100010001001000101010001000100010001000100010001010111100110101010101010101010101010101010101010101011101010111011100101010101010101010101010101010101010101100110011101111000100010011010101010101010101010101011101110111100101110111011101110111011110011001100110010111011101110111011101110100101001101010101001100110010000100010010001000100010001000100001000100010001001000100010001000100010001100110011001100110100010101010110011001110111011101111000100010001000100010000111011101110111011101110111011101110110011001100101010000110100,
	2400'b010101010100010001010110011101110111011101110111011101100111011101110111011101110111011101110111011101110111011001110111011101010010001000100010001101111000100010001000100010011001100110101010101010011001100110101010101010101001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000011001100101010001000100010110001001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001110110011001110110010001000110011101010110011001100111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011101111001100101110111011101111001101110111001011101110111011101110111011101111001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101110111011101101110111011101110111011101110111001100110011001100110011001100110010111011101001100011001100110100010001000100010001000100010001000100001101000110011001100110100010000111011001100101010101000011001000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000010010010001010101010000110100100010000111100001110111011101100110011001010101010101000101010001000100001100110010001000100010001000100010001000100011011001100100010001000100010001000101011110011010101010101010101010101010101010101010101010101001011001010101010101010101010101010101010101100111100010001001100110011010101010101010101010111011101111001100110010111011101110111100110011001100110010111011101110111011101110100101001101010100001100100010001000100010001000100010001000100010000100010001001000100010001000100010001100110011001101000100010101110111011101111000100010001000100010001000100010001000100010001000011101110111011101110110011001100101010001000100,
	2400'b010101010100010101010110011101110111011101110111011101110110011101110111011101110111011101110111011101110111011001110110011101000010001000100010010010000111100010001000100110011001100110101010100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001111000011001100110010101000100010101111001100110011001100010001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001110110011001100101001100110101010101010101011001100111011110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101111001100110010111011110011011101110111011101110011001011101110111011110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101110111011101101110111011101110111011101110111011100110011001100110011001100101110111010011000110011001100110100010101000100010001000100010001000100010001010110011110000111011110011001100010000110010000110010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000010010001101000101010101000011010110001000100010001000100001110110011001010101010101010101010101000100001100110011001000100010001000100010001000100010010001010101010001000100010001000100010101111001101010101010101010101010101010101010101010101000010101010101010101010101010101010101011001111000100110011001101010101010101010101010101110111011110011001100110010111011101110111100110011001100110010111011101110111011101110010100001101010011001000100010001000100010001000100010001000100010000100010001001000100010001000100011001100110100010001010101010101110111011110001000100010001000100010001000100010001000100010000111011101110111011101100110011001100101010001000101,
	2400'b010101010101010101010110011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101100110011000110010001000100011011010001000100010001001100110011001100110011001100110001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000011001100110010101000101010101111000100110011001100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100001110110011001110110010000110100001101000101010101100111100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101111001100110011001100110111011110111011101110111011011101110011001100110111101110111011101110111011101110111011101110111011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110011011100110011001100110011001100110010100110001100110011001101000101010001000100010001000100010001000100010101100111100010011001100110011001100110010110001100100010001100110011001000100010001000100010001000100001000100100010001000100010001000100010001000100010001000010001001000110101011001010011001001101000100110011000100010000111011101100110010101010110011001010101010001000011001100110011001000100010001000100010001000110101010101010101010101010101010101010111100110101010101010101010101010101010101010010110010101010101010101010101010101010110011110001000100110101010101010101010101010101010101110111100110011001100110010111011101110111100110011001100101110111011101110111011101110010100010001010011001000100010001000100010001000100010001000100010000100010010001000100010001000110011001100110100010101010110011001110111100010001000100010001000100010001000100010001000100001110111011101110111011101100110011101100101010001010101,
	2400'b010101010101010101010110011101110111011101110111011101110111011101100111011101100111011101110111011101110111011101100111010100100010001000110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000011101100111010101010101010101111000100110011001100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100001110110010101010111010000110011001100110100010001010111011110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101111001100110011001101110111011110110111101110111011101110110111011110111011101110111011101110111011101110111011101101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011100110011001100110011001100101001100011001100110011001101000101010001000100010001000100010101010101010101111000100010011010101110101010100101110100001100110011001100100010001000100010001000100010001000100001000100100010001000100010001000100010001000100010001000100001001000100011010101100100001000110111100110011000100110001000011101110110011001100110011001100101010001000100010001000011001100100010001000100010001000100011010101010101010101010110011001100101011110011010101010011001100110011001101010000101010101100101010101010101010101100111100010001001101010101010101010101010101010101011101110111100110011001100110010111011101110111100110011001100101110101010101110111011101110010100010001000010001100100010001000100010001000100010001100110010000100010010001000100011001000110011001100110011010101010110011001100111011110001000100010001000100010001000100010001000100001110111011101110111011001110111011101100100010101010101,
	2400'b010101010101010101100110011101110111011101110111011101110111011101100111011101100111011101110111011101110110011001100110010000100010001000110101100010001000100010001001100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101111000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100111010101010110011001111000100110001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000111011101110111011101100101010001000101010000100010001000110011001101000101011110001000100010011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101111001100110011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110011001100110011001001010100110011001100110011010001010101010001000100010001010101010101010110011101111000100110011010101010111010011101000011001100110011001000100010001000100010001000100010001000010001000100100010001000100010001000100010001000100010001000100010001000010010010001010101001100100100100010011001100110001000100001110111011101100110011101110101010101010101010001000011001100110011001000100010001000100011001101000101010101010110011001110110011001111001100110011001100110011001100101110101011001100101010101100110011001110111100010011010101110111010101010101010101010111011101110111011110011001100110010111011101110111100110011001100101110101010101110111011101110000100010000110010001000100010001000100010001000100010001101000010000100010010001000100011001000100011001100110011010001100101011001110111011101111000100010001000100010001000100010001000100001110111011101110110011101110111011101010101011001100110,
	2400'b010101010101010101100110011101110111011101110111011101110111011101100111011001100110011001110111011001110110011001100110001100100010001000110101100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011001010110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010011000100010011001100110011001100110011001100110011001100110011001100110011001100010000111011101100101011001010100001100110011001100100010001000100011001101000110100010000111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101111001100110011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111001100110010010101001100110011001100110011010101010101010001000101010101010101011001110110011110001001101010101001101010101000010000110011001100110010001000100010001000100010001000100010001000010001000100100010001000100010001000100010000100100010001000100010001000100010001000110101010000110011011010011001100110001000100010001000011101110111011101110110011001100101010001000100010001000011001000100010001000100011001100110101010101010101011001100111011001100111100110011001100110011001100101100101011001100101011001100110011110001001101010101011101110111011101010101010101010111011101110111011101110111011101110111011101110111011110011001100101110111011101110111011101101110100010100110010001000100010001000100010001000110011010001000011000100100010001000100011001100110011010001000100010001100110011001110111100010001000100010001000100010001000100010001000100010000111011101110111011101110111011001010110011001100110,
	2400'b010101100101010101100110011101110111011101110111011101110111011101100110011001100110011001110111011001110110011001100101001000100010001000110110100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011000100010001000011101100101010101010100001100110011001100100010001000100011001101000110011101100111100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101110111100110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011001101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011100110011001100100101010011001100110011001100110100010101010101010101010110010101100110011110001000100010011001101010101001100001100100010000110011001100100010001000100010001000100010001000100011001000010001000100010010001000100010001000100010001000100010001000100010001000100010001000100100010100110011010001111001100110011001100010011000100010001000100010000111011101100110010001000100010001000100001100100010001000100011001100110100010101010101011001100111011101110111100010011001100110011001100001010101011101100110011101110111100010011010101110111011101110111011101010101010101010111011101110111011101110111011101110111011101110111011110011001100101110111011101110111011101001100100010000100010001000100010001000100010001100110100010001010011001000100010001000100011001100110011010001000100010001010111011101100111100010001000100010001000100010001000100010001000100010000111011101110111011101110110010101100110011001100110,
	2400'b010101010101011001100110011001100110011101110111011101110110011001100110011001100110011001100111011001100110011001100100001000100010001101000111100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100001110111011101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010011001100110001000100010000111011001100101010001000011001100110010001100100010001000100011001101000110011001100111011110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101110111100110011011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011100110011001001010100110011001100110011001101000110011001010101010101010111011001110111100010011001100110101010101010101001011101010100010000110011001000100010001000100010001000100010001100110011001000010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010010001000011001101101001101010011001100110011001100110001000100110000111011101110111010101000101010101010100010000110010001000100011001101000100010101010101010101100110011101110111011110001000100110011001011101010110100001100110100010011001101010101011101110111011101110111011101010101010101110111011101110111011101110111011101110111011101110111011110010111100101110111011101110111011101001100101001100100010001000100010001000100010001100110100010101000010001000100010001000100011001100110011010001000100010001010111011101110111011110001000100010001000100010001000100010001000100010000111011101110111011101100110011001100110011001100110,
	2400'b010101100110011001100110011001100110011001110110011001100110011001100110011001100110011001100111011001100110011001100011001000100010001101011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000011110001000100001110111011101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111100010001000100001110111011001010101010000110011001100100011001100100010001000100011001101010101010101100111011110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101011101110111011110011011101110111101110111011101110111011101110111011101110111011101110111011011101110111101101110111001011101110111100110011011101110111011110111011101110111011101110111011101110111011101110110111011101111011101110110111011101110111011101110111011101110111011101110010000100001100110011001100110011001101000111011101100110011001101000100010001000100110101001101010111010100110011000011001000100010000110010001000100010001000100010001000100011001100110011001000100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001101000011001101001000100110011010100110011001100110011001100110000111100010000111011001010110011001100100010000110010001000100011010001000100010101100110010101100110011001110111011101111000100010011000011001010111100001111000101010101010101110111011101110111011101110111011101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101001010100001100100011001100100010001000100011001100110100010000110010001000100010001000100011001100110100010001000101010101010111011101110111011110001000100010001000100010001000100010001000100010001000011101110111011101100111011101110110011001100110,
	2400'b011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100011001000100010001101101000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010000111100010001000100010000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001010110011001010101010101100111011101110110010101000100001100110011001000100010001000100010001000100011001101000101010101100111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101110111011101110111011110011001101110111101110111011101110111011101110111011101110111011101101110111001100110111011100110010111011101110111011101111001100110111011110111011101110111011101110111011101110111011101110110111001101110111101101110111011101110111011101110111011101110111011011011101000011001100110011001100110100010001101000011101100110011101111000100110011001101010101001101010111010101001110110010101000101010000100010001000100010001000100011001100110100010001000011001000100001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001101000111100110101010100110011001100110011001100110000111100010001000011101100110011001100101010101000011001000100011010001000100010101100110011001100110011001100111011101110111100010011000010101101000100010001010101110111010101110111011101110111011101110111010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100101010100001000100010001000100010001000100011001101000100010000110010001000100010001000100011001100110100010001010101010101010111011110001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010010001000100010001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010000111011101110111011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100111011101110111011001010101010001000101011001110101010001000100001100110011001000100010001000100010001000100011001101000101010101100111100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101011110011001100110011001100110011001101110111011110111011101110111011101110111011101110111011011100101110111100110010111011101110101010101010101011101110111100110011011101111011101110111011101110111011101110111011101101110011001100110111011101110111011101110111011101110111011101110111000111010001000011001100110011010001000101010101111000011101110111100010001001101010101010101010111010101010111010101010000101010101010100001100100010001000100011001100110011001101000101010101000011001000100001000100100010001000100011001100110010001000100010001100110011001100100010001000100010001000100010001001000110100110101010100110011001100110001001100101110111100010011001100001110111011101110110010101010011001000110011010001010101010101100111011101100110011001100110011101111000100010010111010101111001100110101011110010111011101110111011101110111011101110111010101010101011101110101010101110111011101110111011101110111011101010101011101110111011101110111011101110111011100001010011001000100011001000100010001000100011010001000100010001000010001000100010001000100011001101000100010001010101010101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000010001000100010010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110011001010101010101010101010101100101010101000100001100110011001000100010001000100010001000110011001101000100011001100111100001110111100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101110111100110011001100110011001100110011001101110111101110111011101110111011101110111011101110110111001011101110111011101110111010101010101010101010101010101110111011110011001101110111011110111011101110111011101110110111011100110011001100110011011101110111011101110111011101110111011101101101110101010001000011010001000100010001010110011010001001011101110111100010011001101110111010101110111011101110111011101110000100001101000011001000100010001000100011001100110011010001010110011001010011001000100010000100100010001000110100001100110011001100100011001100110011001100110011001100110010001000100010001000110101100010011001100110011001100110011001100001111000100110011001100001111000100010000111011001100100001100110011010001100110011001100111011101110110011001100110011101110111100001110110011010001010101010111011110010111011101111001011101110111011101110101010101010101011101010101010101010111011101110111011101110111010101010101010101010111011101110111010101010101010011101010011001000100011001000100010001000110011010001010100010101010100001100100010001000100011010001000100010001010101010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110010001000100011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011001100101011001100101010101010110011001010100001100110010001000100010001000100010001000110011010001000101011001110111011101111000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011110011011101110111011100110011001101110111011101110111101110111011101110111011101110111011011101110010111011101110111011101010101010101010101010101010101010101010111011101111001100110111011101110111011101110111011101110111001011101110111011110011001101110111011101110111011101110111011011011001000100010000110100010001000101010101110111011110011001100010001000100110101010101111001011101110111011101110111011101110000011001100110010001000100010001000100011001100110100010101100111011001010011001000100011001000010001001000110100010000110100001100110011001101000011001100110011001100110010001000100010001000100100011110011001100110011010100110011001100110001000100110011001100110001000100010001000011101110110001100110011010001010111011101100111011101110111011101110111011101110111011101100101100010011001101010111011110011001100110010111011101110111011101110101010101010111011101010101010101010101011101110111011101110111010101010101010101110101010101010101010101010101000011001010010001000100011001000100010001000110100010101100101010001010110010000100001000100100011010001000100010101010101011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100010001000100011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110011001100101010101010101010101000011001100110010001000100010001000100010001000110011010001010101011001110110011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011110111011101110111011100110011011101110111011101110111101110111011101110111011101110110111001011101110111011101110101010101010101010101010011010101010101010101010101011101110111011110011001100110011001011110011001100110010111011101110111011101111001100110111001100110111011101110111000111010001000100001101000100010001100111011001111000011110011001100110011001101010101011101111001100110011001100110010111011101110000100001100100010001000100010001000110011001100110100011001110111011001010011001000100010001000100010001000110100010001000100010001000100010001000100010000110011001100110011001100100010001000100100011110011001100110011010101010101010100110001000100110011001100110001000100010011000100010000111010100110100010001010111100010000111011101110111011101110111011110000111011101100110100110011001101010101011101111001100110011001011101110111011101110111010101110111010101010101010101010111011101110111011101110101010101110111011101110101010101010101001100110010110011001000010001000110011001000100010001000110100010101100110010001010101001100100001001000100011010001010101010101010101011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000100010001000110100011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001111000011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100110011001010100010001000011001100110010001000100010001000100010001000110011010001010110011001010111011110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101100110111011101110111011101110111011101110111011101111011101110111011101110111011101101110111001011101010101010101010101010100110011001100110011001100110011010101010101010101110111010101110111010101010101010101010111011101110101010101010101011101110111100110011001100110011011101110010000100010101010100010001000100010101110111011010001000100010101001100110011010101110111011110011001100110011001100110011001011101110010100001100100010001000100010001000110011010001000101011101110111011101010011001000010001000100010010001101000101010101010101010101010101010101000100010001000100001100110011001100110010001000100011011010001010101010101010101010101010101010011001101010011001100110011001100110011000100010011000011101000100010001000110100110011000011101111000011101110111011110000111011101100111101010101001101010101011101111001100110011001011101110111011101110111011101110101010101010101010101010101011101110111011101110101011101110111011101010101001100110011001100110000101011000110010001000110011001100110011001100110101011001100111011001100110010000100001000100100011010101010101010101010101011001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100100010001000110101011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100111011001100100010000110011001100110010001000100010001000100010001000110011010001100101010101100111011110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010111100110111011101110111011101110111011101110111101110110111011101110111101110111011101101110111001010101010101010101010011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011110011001100110011011101101001010101011001000100010001010101011010000111011110001000100110101010101010101010101111001100110011011100110011001100110011001011101110100100001000100010001000100010001000110011010001010110011110001000011101010011001000010001000100010010001101000101011001100110011101100101010101010101010001000100010001000011001100110010001000100010011010001001100110011010101010101010101010011001101010011001100110011001100110011001100110011001100001100101010101000101011110011001100001111000100001111000100010001000011101101000101110111010101010111011101110111100110011001100101110111011101110111011101110101010101010101010101010101011101110111011101010101010101110101010101010011001100110011001100101110110010100110010001000110011001100110011010001000101011001100111011101110111010000100001000100100011010101010101010101010110011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000110101011101100111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100110011001100100001100110011001100110010001000100010001000100010001000110100010101000100010101010110011001111000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010111100110111011101110111001100110111011101110111011101110111011101110111101110110111011101110010111010101010101001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101011101111001100110011011100011101010110011001010101010101010101011110010111100010011000100110101010101010101011110011001101110111011100110011001100110011001100101110010100001000100010001000100010001000110011010001100111100010001000011101100100001000010001000100010010010001100110011101110111011101110101011001100110010101010101010001000100001100110011001000100010010110011001100110101010101010101010101010101010101010011001100110011001100110011001100110011001100110010111011101010101011010011001100110001000100010001000100010011001100001111001101110111011101110111011101110111100110011001100110010111011101110111011101010101010101010101010101010101010101110111011101010101010101010011001100110011001100110011001100001100110010100100010001000110011001100110100010001010101011001110111011101110111010000100001000100100010010101100101010101100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000010010001000110110011101100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011001010011001100110011001100110011001000100010001000100010001000110100010001000100001101000100010101100110011101110111011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011110011001100110011001100110011001101110111011101110111011101110111011101110111011100101110111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101110111100110011001001011001100111011001100110011001100110100010010111100010011001100110101010101010111011110011001101110111011101110011011100110011001100101110000011001000100010001000100010001000110100010101111000100010001000100001100101001000010001000100100011010101100111100010001000100001110110011101110110011001100101010101010100010000110011001000100010010010001001100110101010101010101010101010101010101010011001100110011001100110011001100110011010101010011000100001100101010110001001101010001000100010001000100110011010100001111010101110111011101110111011101111001100110011001100101110111011101110111011101010101010101010101010101010101010101010111010101010011001100110011001100110011001100110001000100001100110010000100010001000110011001101000100010101010110011001110111011101110111010000100001000100010010010001100110010101100110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100011000100100010001001000110011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100001111000011101111000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011001000011001100110011001100110011001000100010001000100010001000100011001100110011001100110100010001010110011001111000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011101110111100101110111011110011001101110111101110110111011101110111011100110010111011101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010111011101110110111011001100111011001110110011001100110100010011000100110101001101010101010101110111011110011001100110111011100110011011100110011001100101001010010001000100010001000100010001100110100011110001001100010011001100001110110001100010001001000100100011001111000100010001000100010000111100001110111011101110110011001010101010001000100001100100010001001111000100110011010101010101010101010101011101010011001100110011001100110101001101010101010101010101001100101110110010101101001101010010111100010011001101010101010100110011010101111001011110010111011101111001100110011001011101110111011101110111011101010101010101010101010101010101010101010101010101010011001100110011001100110011000100010001000100001110110001100100010001100110011001101000101010101100110011101110111011101110111010000100001000100100010010001100110010101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001101000111011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100001111000011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011001000011001100110011001100100011001000100010001000100010001000100010001000100011001100110100010001010110011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010111011101110111011101111001100110111101110111011011101110011001011101110111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101011101110100111011101111000011101110111011001110111100110011000100110101010101010101011101110111011110011001100110111001101110111001100110011001100011100110010001000100010001000100010001000110110100010011001100110011001100110000111001100010001000100100101100010001001100110011001100110001000100010001000011101110111011001100110010101000100001100100010001001011000100110011001100110101010101010111011101010011001100110011001100110101010101010101010101010101001100110010111011001101000101010011000100010101010101010111011101010011011101111001100110011001011101111001100110010111011101110111011101110111011101110101010101010101010101010101010101010101010100110011001100110011001100110001000100010001000100010000101001100100011001100110011001101000101011001100110011101110111011101110111010100110001000100100010010001100110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010010000100100010001101010111011001100110011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110101010101010100001100110011001100110011001000100010001000100010001000100010001000100011001101000101011001110111100010001000100010001000100110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101011101110111100110111101110111011011100110010111011101110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010010111100010001000011110000111011101110111100110011001101010101010101010101010101110111011101111001100110011001101110111011100110011001010010000100010001000100010001000100010001101001000100110011001100110101010100110010111001000010001001001000111100110011001100110011001100110011001100110001000100010001000011101110110010101100100001100100010001000111000100110011001100110101010101010111011101010011001100110011010101010101010101010101010101010101010100110011000011101101000100110101000100010101010101110111011101010101011110011001100110011001011110011001100101110111010101010101010101010111011101110111010101010101010101010101010101010011001100110011001100110011001100010001000100010001000100001110100001000100011001100110011010001000101011001100111011101110111011101110111011101010001000100100011010001100111011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000010000100100010010001100111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100001111000100001110111011101110110010101010100010001000100010001000011001100100010001000100010001000100010001000110011010001010110011101110111100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101110111100110111101110110111011100101110111011101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010001000100010001000100010000111100010001000100110011001101010101010101010101010101010111011101110111011110011001101110111011100110011000111001000100010001000100010001000100010001101101001100110101010100110101010101010010110001000010001001101101000100110011001100110011001100110011001100110011000100110001000100001110110011001100101001100100010001000100110100110011001100110101010101010111011101010011001100110101010101010101010101010101010101010101010101010011000100001111000101010101001100110101011101110111011101110111011110011001100110011001100110011001100101110101010101010101010101010101011101110111010101010101010101010101001100110011001100110011000100010001000100010001000100010001000100001110011001000110011001100110100010001010101011001110111011101110111011101110111011101100010000100010011010001010111011001100111011110001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110010001000100011010001110111011001110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110010101010101010001000100010001010101010001000011001100100010001000100010001100110010001100110100010001010101011001100110011101110111011101110111100010001000100010001000100010001001100110011001100110011001100110011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010111011110011011101110111001011101110111010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001100010001000100010001000100110011001101010101010101010101010101010101010101010101011101111001100110011001100110010000011001000100010001000100010001000100011010001111001101010101010101010101010101010010101000100010001010101111001100110011001100110011001100110011001100110011001100110011001100010000111011101100101001100110010001000100011100010011001100110101010101010111010100110011001101010101010101010101010101010101010101010101010101010101001100001111000101010101001100110101011101110111011101110111011101111001100110011001100110011001011101110101010101010101010101010101011101110111010101010101010101010101001100110011001100110011000100010001000100010001000100010001000011101010011001100110011001100110100010001010101011001110111011101110111011101110111011101100010000100100011010001010111011001100111100010001000011101110111011101110111011110001000011110001000100010001000100010001000100010001000100010000111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100110011010000110011010101110111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010000111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001110111011101100101010101000100001101000100010001000100010001000100010001000011001000100010001000100010001100110011010001000101010101010101011001100110011101110111011101110111100010001000100010001000100110011001100110011001100110011001100110011001100010000111100110011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101011101111001100110010111011101110111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100010011000100010011001101010101010101010101010101010101010101010101010101010101010101110111100110011001100100101000010001000100010001000100010001000100011010101111010101010101010101010101010101010010100000100010010011010001001100110011001100110011001100110011001100110011001100110011001100110011000011101110100010000110011001000100010010010001001100110011010101010101010100110011001101010101010101010101010100110101010101010101010101010101001100110001000101010101010101010101010101010111011101110111011101110111100110011001100101110111011101110101010101010101010101010101010101110111010101010101010101010101001100110011001100110001000100010001000100010001000100010000111011001000011001100110011001100110100010101010101011001110111011101110111011101110111011101100010000100100010010001010111011101110111100010001000100001110111011101110111100010001000100001111000100010001000100010001000100010001000011101110111100010001000100010001001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000110100010101000100011001110110011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001010101010001000100010001000101010101010101010101010101010101000011001100100010001000100010001000100011010001010101011001100110011001110111100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110001000100001110111100010011001100010001000100010001000100110011001100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101110111011101110111011101110111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011000100110011001100110101010101010101010101010101010101010101010101010101010101010111011101110111010010100110010001000100010001000100010001000100011010101111001101010101010101010101010101010000011000100010010011010001001100110011001100110011001100110011001100110011001100110011001100110011000100001100101010101000011001000100010001001011000100110101010101010101010100110011010101010101010101010101010101010101010101010101010101010101010100110001001101010101010101010101010101010101010101010111011101110111011101110111011101110111011101010101010101010011001100110101010101010101010100110011010101010101001100110011001100110001000100010001000100010001000100001110110010100110011001100110011001100110100010101010110011001110111011101110111011101110111011101110010000100100010010101010111100010001000100010001000011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100110011010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000110100010101000101011101110111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100110010101010101011001010110011001100110011001010100001100110011001000100010001000100010001000100010001100110100011001100101010101100111011110001000100010001000100010001000100010001000100010001000100110011001100110011001100010001000011101100110011110001001100001111000100010001001100110011001100110011001100110001001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101110111011101110111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101110100110001100110010001000100010001000100010001000110011010110001001101010101010101010101010101010000010000100010010010110001001100110011001100110011001100110011001100110011001100110011001100110011000011101010111010101000011001000100010001000110111100110011001101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010101010101010101011101110111011101010101010101010101010100110011001100110011010101010011001100110101010101010101001100110011001100110001000100010001000100010001000100001110111010100110011001100110011001101000100010101010110011001110111011101110111011101110111011101110010000100100010010101100111100010001000100010001000011101110111011101110111011101111000100010001000100001111000100010001000100010001000100010001000100010001001100110011010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100001000100011010001000110011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010000111100001111000100001111000011110001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100110011001100110011001100110011001100110010101000011001100110011001000100010001000100010001000100010001000100011010001010110011001100110011110001000100010001000100010001000100010001000100010001000100010011001100110011000100010000111011101100110011010001000011101100110011010001000100001110111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101011101110111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010100101100100001100110010001000100010001000110011001100110011010010001001100110101010101010101010101001110010000100010010011110011001100110011001100110011001100110011001100110011001100110011001100110010111011001110111010101000100001100100010001000110101100010011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001100110011001100110011010101010101001100110011001100010001000100010001000100010001000100010000110010000110011001100110011001101000101010101100110011101110111011101110111011101110111011101110011000100100010010101100111100010001000100010001000100010001000011101110111011110001000100010001000100010000111100001111000100010001000100010001000100110011001100110101010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100011001000100010001101010110011101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010000111100010001000011110000111100010001000100010001000100010001000100010000111100010001000100010000111011101110111011101110111011001100110011001100110011001100100001100110011001100110011001000100010001000100010001000100011001100100010001100110100011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001010101010101111000011101010101010101100101010101010110011001111000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101110111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101001011101000100001100110010001000100010001100110011001101000100001101111001100110101010101010101010101001100010000100010011100010011001100110011001100110011001100110011001100110011001100110011001100110000110011110000110010101010100001100100010001000110011011010011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100001110101010000110011001100110011001101000101011001100110011101110111011101110111011101110111011101110011000100100010010101100111011110001000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110101010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000100100010001101010110011101110111011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010000111100001111000011110000111011110001000100010001000100010001000100010001000100001111000100010000111011101110111011101110111011101100110011001100110011001000011001100110011010001000011001000100010001000100010001000100011010000110011001100110011010001010111011110001000100010001000100010001000100010001000100010001000011110001000100010001000100010000111011001010101010101010111011001010100010000110011001101010110011010001000100010001000100010001000100110001000100010001001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101011101110111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110010111010101010100001100110010001000100010001100110011001101000101010001011001100110101010101010101010101001010001000100010100100110011001100110011001100110011001100110011001100110011001100110011001100001111000100110000110011001100101001100100010001000110011010110001001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110101001101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100001110101001100110011001100110011010001000101011001100110011101110111011101110111011101110111011101110100000100100011010101110111011101111000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010010000100100011010001010111011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000100010000111011101110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110110010000110011001100110011010001000011001000100010001000100010001000100011010001000011001100110011001100110101011001111000100010001000100010001000100010001000100010001000100001110111100010001000100001110110010101010101010101010110011001010100001100110011010001010101011110001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010111011110010111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110011010100110011001100110000111011001010100001100100010001000100011001100110011001101000101010101011000101010101010101010101010100101010001000100010101100110011001100110011001100110011001100110011001100110011001100110011001100010001001100101110111011001100101010000100010001000110011010001111001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100001110100001100110011001100110100010001000110011001110110011101110111011101110111011101110111011101110100001000100011010101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000010001000100010010001100111011001100110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010000111011101110111011110000111011101111000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011001010011001100110011001100110100010101000011001000100010001000100010001000100011001101000100001100110011001100110011010001010111100010001000100010001000100010001000100010001000100010000111011110001000100010000110010001000100010101010101011001000011001100110011010001000101011110001000100010001000100010001000100010001000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101110111100101110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111010101000011001100100010001000100011001100110011001101010110010101010110100110101010101010101010100101000001000100100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001110111011001100110010000100010001000110011001101101000100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100001100100001100110011001101000100010001010110011101110111011101110111011101110111011101110111011101110101001000100011010001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110010000100010010010001100111011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011110001000100001110111011101111000011101110111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110010000110011001100110011001100110100010000110010001000100010001000100010001000100011001101000101010000110011001100110011010001000101011010001000100010001000100010001000100010001000100010001000011001100111100010000110010101000100010001000100010000110011001000110011001101000110011110001000100010001000100010001000100010001000100010001000100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011101111001100101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110010110010100110011001100100010001000100011001101000100010001000111011001100110011110101010101010101010100100110001000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110000111011001110110010000100011001100110011001101011000100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000011101010100001100110011010001000100010001010110011101110111011101110111011101110111011101110111011101110100001000100010010001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001000100100011010101100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111100010000111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100001110111011101110111011101100100001100110011001101000011001101000100010000110011001000100010001000110011001000100011001100110101010101000011001100110100010001000100010101101000100010001000100010001000100010001000100010001000011101100101011101110110010101000100001100110011001100110011001100110011001101000110011001110111100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011110011001011101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000101010000110011001100100010001000100011010001000100010001000111100001100111011110011010101010101010100000110001000100111000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000111011101110110010000110011001100110011001101000111100110011001100110011001101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001001100110011001100110011000100010001000100010001000100010001000100010001000100010001000011101010100001100110100010001000100010001010110011101110111011101110111011101110111011101110111011101110011001000100010001101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100010001000110100010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000100010001000100010001000100010001000100010000111011101110111011001000011001100110011010001000100010000110100001100110011001000100010001000110011001000110011001100110100010101010100001100110100010001000100010101100111100010001000100010001000100010001000100010001000100001110110010101100110010101000011001100110011001100100010001000110011010001010110011001111000100010001000100010001000100010001000100010001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101100110011001010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100100001100110011001100100010001000100011010001000101010101000110100110000111100010001010101010101010100000110001000101001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110010111011101110110010000110011001100110011001101000110100010011001100110011010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010001000100010001000011101010100001100110100010001000100010001100111011101110111011101110111011101110111011101110111011101110100001000010010001101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000100010001001000101011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110110011001110111011110001000100010001000100010001000100010001000100001111000100010000111011101110110010000110011001101000100010001000100010001000100001100110011001000100010001000110011001000110011001100110100010101100101010001000100010001000100010101010110100010001000100010001000100010001000100010001000100010000111011001010100010000110011001100110011001100100010001000110011010001010110011101111000100010001000100010001000100010001001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010111100110010111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001010100001100110011001100110010001000100011010001010110011001100110100110010111100110101010101010101010011100100001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001110110001101000100010000110011001101000101100010011001100110011001100110011010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100010000111010101000100010001000100010001010101010101100111011101110111011101110111011101110111011101110111011101110100001000010010001101100111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000100010001101010101011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011101110111011101100110011001110111011101110111100010001000100010001000100010001000100010001000100001110111011101100100001100110011010001000100010001000100010001000100001100110011001000100010001000110011001000110011001100110100010101100110010101000100010001000101010101100110011110001000100010001000100010001000100010001000100010001000100001110101010000110011001100110011001100110010001000110100010101010110011001110111100010001000100010001000100010001000011101111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101000011001100110011001100110010001000100011010001010110011110000111100010101001100010101010101010101010011100100001001001101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001110101001101010101010000110011001101000101011110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100010001000100010001000100010000111010101000100010001000100010001010101010101100111011101110111011101110111011101110111011101110111011101110101001000010001001001100111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100100011010101010110011001100110011001100110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010111011101110111011001100111011001010110010101100111011101100110011110001000100010001000100001110111011110001000100001110111011001000011001100110100010001000100010001010101010101000100001100110011001100100010001001000011001000110011001100110100010001100110011001010100010001000101010101100111011110001000100010001000100010001000100010001000100010001000100010000111010100110011001100110010001000100010001000110100010001000100010101100111011101110111011110001000011101100110011001111000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010101000011001100110011001100110011001000100011010001010111100010001000100010101001100110101010101010101001011000100001001001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000100010101100101010101000011001101010110011110001001100110011001100110011001100110101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010000110010101000100010001000100010101010101011001100111011101110111011101110111011101110111011101110111011101110101001000010001001001010111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000100011010101100110011001100110011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101000100011001110111011001010101011001010101010101010110011001010101011101111000100010001000011101110111011110001000100001110110010000110011001100110100010001000101010101010101010101000100010001000011001100100010001000110011001100110011001101000100010001100110011001010101010001010101010101100111011110001000100010001000100010001000100010001000100010001000100010000111010101000011001100100010001000100010001100110100001100110100010101100111011101110111011101110110011001100110011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110010000110011001100110011001100110011001100110011010001010111100010001001100110101010101010101010101010101001011000100001001001111001100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110001000100001110100011101110101010101000100001101010110011010001000100010011001100110011001100110101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110001000100010001000100010001000100010001000100010000111010101000100010001000100010101100101011001100111011101110111011101110111011101110111011101110111011101110110001000010001001001010111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100100001000100011010101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101000100010001010110011001100100010001000100010001010110011001000101011001110111011101110111011101110111011110000111011101110101010001000100010001000100010101010101010101100110010101010100010101010011001100100010001000100010001100110011001101000100010001010110011101100110010101010101011001100111100010001000100010001000100010001000100010001000100010001000100010000110010000110011001000100010001000100010001000100011001100110100010101100111011001100110011001100110011001100111011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000101010000110011001100110011001101000011001100110100010101010111100110011001100110101010101010101010101010101001010100100001001110001001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011000100001110110100001110110010101000011010001010111011101111000100010011001100110011001100110011001101010101010101010101010101010101010101010101010100110011001100110011001100110011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000100010001000100010001000100010001000100010000111010101000101010001010100010101100101011001110111011101110111011101110111011101110111011101110111011101110110001000010001001001010111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100100001000100011010101100111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101000100010001000100010101010101010000110100010001000101010101000101011001100110011001110111011101110111011001100110011101110110011001010100010001000101010101010110011001100110011001010101010101010011001000100010001000100010001000110011001101000100010001010110011101110110011001010101011001100111100010001000100010001000100010001000011101110111011101110111011101110100001100110010001000100010001000100010001000100010001100110101011001100110011001100110011001100110011001110111011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001100101010101000011001100110100010001000100001100110100011001100111100110011001101010101010101010101010101010101001010100100001001110001001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001100001100111100001110110010100110011010001010111011101111000100010001000100110011001100110011001101010101010101010101010101010101010101010101010100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000100010001000100010001000100010001000100010000111010101010101010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111001000010001001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001010011001000110100010101100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101000100010001000100010001000100001100110011001100110100010001000101010101010110011101110111011101110110010101010101011001110110010101000100010101010101011001100110011001110111011001100110011001000011001000100010001000110011001100110011001101000100010001000110011101110110011001100101011001111000100010001000100010001000100001110110011001010101010001000100010001000101010000110010001000100010001000100010001000100010001101000101010101100101010101100110011001100110011001110111100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101100110011001000011010001000100010001010101010001000101011001110111100110011001101010101010101010101010101010101001010000100001010010011001100110011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100001111000100001110110010100110011001101010111011110001000100010001000100110011001100110011001101010101010101010101010101010101010101010101010100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110001000100010001000100010001000100010001000100010000111010101010101010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111001100010001000101000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001010010001000110100010101100110011001100110011001100110011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010001000100010001000101010000110011001100110010001000110011001100110100010001010110011101110111011001010100010001010110011001100101010101010101010101010110011001100110011001110111011001100110011001000011001100100010001100110011001100110011001101000100010101010101011101110111011001110110011001111000100010001000100010000111011101100110010101010101010001000011001100110011001100110011001000100010001000100010001000100011010001010101010001000100010001010110011001100110011101110111100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101110111010101000011010001010100010101100110011001100110011101111000100110011001101010101010101010011001100110101000010000100001010010011001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001011110001000100001110110010100110011001101010111100010001000100010001000100010011001100110011001101010101010101010101010101010101010101010101001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110001000100010001000100010001000100010001000100010000111010101010110010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111001100010001000100110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001000010001000110100010101100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010100010001000100010001000100010101000011001100100010001000100010001000110011010001010110011101110110010101000100010101100110011001100110011001100110010101100110011001100110011101110111011001110111010101000011001100110011001101000011001100110011010001000101010101010101011101110111011101110110011001111000100010001000100001110111011001100110011001100110011001000100001100110010001000100011001100100010001000100010001000110011010001010100001100110100010001010110011001100110011101110111100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101110110010001000100010101010110010101101000011101110111011110001000100110011001100110011001100110011001100110101000001100100001010110011001100110011001100110101010101010101001100110011001100110011001100110011001100110011001100110011001100010011001011101110110010100110011001101010110100010001000100010001000100010001001100110011001100110011001101010101010101010101010101010011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010000111010101100110010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111010000010001000100110110100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011000110010001000100100010101100110011001100110011001100110011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100010000110011001100110011010001010100001100110010001000100010001000110011010001010110011001100101010001000100010101100110011001110111011001100101011001110111011101110110011101110110011101110111010101000011001100110011010001000100001100110100010001000101011001010101011110001000011101110111011001111000100010001000100001110111011001100111100001110111010101000100001100110010001000100010001000100010001000100010001000110100010000110011001100110011010001010110011001100111011101111000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101100101010101000100010101100111011001111000100010001000011110001001100110011001100110011001100110011001100110011000001100100001010110011001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100110011000100010011000011101110110010101000011001101000110011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010000111010101100110011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111010000010001000100100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110010100100010001000100100011001110110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110010101000011001100100010001100110100010000110010001000100010001000110011010001010110011001010100010001010101010101100111011101110110011001100110011001100111011101100110011101110110011101110110010101000011001100110011010001000100010001000100010001010101011001100101011110001000011101110111011001111000100010001000100010000111011101111000100001110110010101000011001100110010001000100010001000100010001000100010001000100011001100100010001100110011010001000100010101100111011110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011001010110010101000100011001100111011101111000100010011000011110011001100110011001100110011001100110011001100110010111001100100001010110011001100110011001100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110000111011101110110011001000011001100110110011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010000111010101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100010001000100100110100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110010100100001001000110101011001100110011001100110011001100110011001100110011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010100110011001100100010001000100011010000110010001000100010001000110011010001010101010101000100010001010101010101100111011101110111011101100110011101110111011001010110011101100110011101110110010101000011001100110100010001010100010001000100010001010110011101110110011010001000100010001000011101111000100010001000100010001000100010001000100001110101010001000011001100110011001000100010001000100010001000100010001000100011001000100010001100110011001101000100010101100111100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110010101010110010101000101011001111000100001111000100110011001100010001001100110011001100110011001100110011001100110010111001100100010011010011001100110011001100110011001100110101001100110011001100110011001100110011001100110011001100110011001100110000110011101111000011001000011001000110110011101111000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100010001000100010001000100010000111010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000010001000100100101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110010000100010001000110101011101100110011001100110011001100110011001110110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010001000011001100100010001000100010001000110011001000100010001000110011010001000100010001000100010001000101011001100111011101110111011101110111011101100110011001100111011101100110011101110110010101000011001100110100010001010101010001000100010001010101011101110111011010001000100010001000011101111000100010001000100010001000100010001000011101100101010101000100001100110010001000100010001000100010001000100010001000100011001000100010001100110011001100110100010101100111100010001000100110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000110010101010110011001010101011001111000100010001000100110011001100010011001100110011001100110011001100110011001100110010111001100100010011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001100111100010001000011000110011001100110101011101110111100010001000100010001000100010001001100110011001100110011001100110011000100010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011000100001000100100101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110001100010010001001000110011101100110011001100110011001100110011001100111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101000100010101000100001100110010001000100010001000100010001000100010001000100011001101000011001100110100010001010101011001100111011101110111011101110111011101110111011001100110011001010101011001100101010001000011001100110100010001010101010001000100010001010101011001110111011010001000100010001000100001111000100010001000100010001000100010001000011101100101010001000100001100100010001000100010001000100010001000100010001000110011001000100011001100110011001100110100010001010101011001110111100010001000011101111000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110110010101100110011001010101011101111000100010011000100110011001100110011001100110011001100110011001100110011001100110010111001100100010011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101111000100010001000011000110011001000110101011110001000100010001000100010001000100010001001100110011001100110011001100010001000100010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101110111011101110111011101110111011101110111100010001000011101110111011101110111011101110111011000100001000100010100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100101001000100001001001000110011101100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101000101010001000101010001000100001100100010001000100010001000100010001000100010001000100010001100110011001100110100010101010110011001100111011101110111011101110111011101110110010101000100010101000101010101000101010001000011001101000101010001010101010101000100010001010101010101100111011010001000100010001000100010001000100010001000100010001000100010001000011101100101010101000011001100100010001000100010001000100011001000100010001000110011001000100011001100110011001100110100010001010110011101110111011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001100110010101100110011001100110011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110010110001100100010011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100110001000011000110011001100110100011110001000100010001000100010001000100010001001100110011001100110011000100010001000100010001001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100001000100010100011110001000100010001000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100100001000010010001101010110011101100110011001110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001000100010000110011001100110011001000100010001000100010001000100010001000100010001000100010001100100011001101000101010101010101010101010110011101110111011101110111011101100100010001000100010001000100010101010101010001000011001101000101010101010101010101010100010101010101010101100111011001111000100010001000100010001000100010001000100010001000100010000111011101100101010101000100001100110011001100100011001100110011001100100010001000100011001100110011001100110011010001000101011001110111011110001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101100110011001100110011001110110011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110010101001000100010011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000011001000011001100110100011110001000100010001000100010001000100010001001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010011011110001000100010001000100010001000100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100011001000100010001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101000100010000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100011001101010101010101010101010101100110011101110111011101110110010101000100010001000100010001000100010101010101010000110011001101000101010101100101010101010101010101010101010101100110011001111000100010001000100010001000100010001000100010001000100010000111011101100110011001010100001100110011001100110100010001000100010000100010001000100011001100110011001101000100010101100111011101111000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011001110110100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110010100001000100010011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000011001000100001100110100011110001000100010001000100010001000100010001000100010001001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011100110001000100010011011110001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100011001000100010010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010001000100010001000011001100100010001000100010001000100010001000100010001000100010001000100010001000100100010001000101010101010101011001100110011101110111011101110101010001000100010001000100010001000101010101010101010001000011010001010101010101100110011001100101010101010101010101100110011001111000100010001000100010001000100010001000100010001000100010000111011101100110011001010101001100110011001100110100010101010101001100100010001000100011001100110100010001010101011001100110011101110111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011110000111100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000100011011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101000100001101000100011110001000100010001000100010001000100010001000100010001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010010011010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001010010001000100010010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010001010100010001000011001100110010001000100010001000100010001000100010001000100010001000100010001000110100010001000101010001000101011001100111011101110111011001100101010101010101010101010101010101010100010101010101010001000100010001010101010101100110011001100101010101010101010101100111011001111000100010001000100010001000100010001000100010001000100010000111011101110111011101100101001100110011001100110101011001100011001000100010001100110011001100110100010001010110011001100110011001110111100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110000011001000100011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101000100001101000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010010011010001000100010001000100010001000100001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001000010000100100010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101010101000100001100100010001000100010001000100010001000100010001000100010001000100010001000110100010001000100010001010110011001100111011101110111011101100110010101010100010001000100010001010100010101010101010001000100010001010101010101100110011101110110011001010101010101100111011110001000100010001000100010001000100010001000100010001000100010001000011101110111011001010100001100110011001101000101011001000010001000100010010101100101011001010100010001010101011001100111011101110111011101111000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100001110111100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110000011001000100011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101010100010001000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101000001000100010010010110001000100010001000100010001000100010000111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011000110001000100100011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100101010101000100001100100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001010110011101100110011001110111011001100100010001000100010001000100010001000101010101010101010001000100010101010101011001100110011101110111011001100110011001100111011110001000100010001000100010001000100010001000100010001000100010001000011101100101010001000011001100110100010001100110010000100010001000100010001101010110011101110110010101010101010101010110011101110111011101110111100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110000011001000010011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101010101010001000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101010001000100010001010101111000100010001000100010001000100010001000011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110010100100001000100100011011010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100101010101000011001100110010001000100010001000100010001000100010001000100010001000100010001101000100010000110100010101010101010101000100010001000101010101010101010001000100010001010101010101010101010101010101010001000100010101100110011001100111011110000111011101100110011001101000100010001000100010001000100010001000100010001000100010001000100010000110010101000100001101000100010001000101011001100100001000100010001000100010001000110100010001000100010001010110010101010101011001111000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110011001000010011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101010110010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101010001000100010001010001111000100010001000100010001000100010001000011101110111011101110111011101111000100010001000100001111000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110010100100001001000100100011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010100110011001100110010001000100010001000100010001000100010001000100010001000100010010001000011001100110011001100110011001101000100010001000100010101010101010101010101010101010101010101010101010101010101010001000100010101100110011001110111100010001000011101110111011001111000100010001000100010001000100010001000100010001000100010001000011101010100010001000100001101000100010001100110011001010011001000100010001000100010001000100011001100110011001100110100010101100101010101010110100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110011001000010011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101100110010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000111011101110111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111100001100010000100010001010001111000100010001000100010001000100010001000100001110111011101110111011101110111100001111000011101111000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110001100010001000100110101011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100100010001000100001100110010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001000100011010001100110010101010101010101010100010101010101010101010101011001100101010101100101010001000100010101100110011001110111100010001000100001110111011001111000100010001000100010001000100010001000100010001000100001110110010001000100010001000100010001000101011001100110010101000010001000100010001000100010001000110011001100110011001100110100010001010110011001010101010101111000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110011001000010100100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100001110110010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111100010000111011110000111100001110111011101110111011101110111011101110111011101110111011101100010000100010001001101111000100001111000100010001000100010001000100010001000011110000111011101110111011101110111100001111000100010001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110001000010001001000110110100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000100010001010100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001100111011101100110010101000100010101010110010101010101010101100110010101100101010001000101010101100110011101111000100010001000100010000111011101111000100010001000100010001000100010001000100010001000011001010100010001000100010001000100010001010111011101100110010100110010001100110010001000100010001000110011001100110011001101000100010001000101011001100110010101010110011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110011001000010100100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100010011000100001110111011001010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001111000100010001000100010001000100010001000100010001000100010000111011110001000100010000111100010001000100010001000100010001000100010000111,
	2400'b011001100110011001100110011001100110011001100110011001100101001000010001001001000110100010000111011101111000100010000111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010000111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010001000101010101010100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001010111011101110111011001010100010001010110011001010101011001100110010101010101010001000101010101100111011101111000100010001000100010000111011110001000100010001000100010001000100010001000100001100101010001000100010001000100010001000101011001100111011101100101001100110011001100100010001000100010001000110011001100110011001101000100010001000101010101100111011001010100010101101000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110010001000010100100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100001110111011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010000111100010000111011101110111011101110111011101110111011101110111011101110111011101110010000100010001001001101000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011110000111100010001000100001111000100010000111,
	2400'b011001100110011001100110011001100110011001100110011001100100000100010001001001010111100010000111100010001000100010001000100010001000100001110111011101110111011101110111011101111000100010001000100010001000100010001000011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010001010110011001010100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011010001010111011101110111011101100101010101010101011001010101011001010110011001010100010001000101010101100111011101111000100010001000100010000111100010001000100010001000100010001000100010000111011001000100010001000100010001000100010001000110011101110111011101100100001100110011001100100010001000100010001000110011001100110011001101000100010001000100010101100110011001100101010001000101100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110010001000010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110011000100010000111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001001001101000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100011000100010001001101101000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011110001000100010001000100010001000100010001000100001110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010100001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010101010111011101110111011101110110011001010100010101010101010101100111011101100100010001000101010101100111011110001000100110011001100110001000100010001001100010001000100010001000100001100110010101000100010001000100010001000101010101100111011101110111011101100011001100110011001000100010001000100010001000110011001100110011010001000100010101000101011001010101010101010110010101010100010101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000010101100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001100110011001100110011000100110001000100010000111011101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001001001010111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001110110011001100110011001010010000100010001010001101000100010001000100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110000111011101111000011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010000110010001000100010001000100010001000100010001000100010001000100010001000100011001100110100010001000101011001100111011101110111011101110111011101100101010001000100010101100111100001100100010001010101010101100111100010001000100110011001100110011000100010001000100010001001100010000111010101010101010101000100010101000101010101000101011001110111011101111000011101000011001100110011001100100010001000100010001000110011001100110100010001000100010101010101010101010101010101010101010101010101010101010111100010011001100110011001100110011001100110011001100110011001101010011001101010101010100110011010101010011010101010011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001000101000111100010000111011110001000100010001000100001111000100010001000011101110111011101110111011101110111100010000111011101110111011101110111,
	2400'b011001100110011001110111011001100111011101100110011001000010000100010010010101111000100010001000100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101000011001000100010001000100010001000100010001000100010001000100010001100110100010001000100010001000100010001010110011101110111011101110111011101110101010001000100010101100111011101010100010001000101011001110111100010001001100110011001100110011001100110001000100110011001100001110101010001010101010101010101010101010101010101010110011101110111011110001000010100110011001100110011001000110010001000100011001100110011001101000100010001010100010101010101010001000100010101010110011001100110011001100110011110011001100110011001100110011001100110011010101010011001100110101001101010101010100110011010101010011010101010101010101010101001100110011001100110011001100110011001100110011001100110101001100110011001100110011001101010101010101010011001101010011001101010101001100110011001100110101010101010101010101010011001100110011001100110101010101010101001100110011001100110101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000101000111100010000111100010001000100010001000100001111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001110111011101110111011101110111011101110111011000110001000100010010010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010001000100010001000011101110111011110001000100001110111011101110111011101100110011001010101010101000100010001000100010001000100010101100110011001010011001100110011001101000011001100100010001000100010001000100010001100110011001100110011001101000100001100110100010101100111011101110111011101110110011001000101011001110111011101010100010001010101011001111000100010011001100110011001100110011001100110011001100110011000011101010100010001010101010101010101010101100101011001100111011101110111011110000111010000110100001100110011001100110011001100110011001100110011001100110100010001000100010101010101010001000100010101010110011001100110011101100110011001111001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001101010101010101010101010101010101010100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000100110111100001111000100010000111100010001000011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011101110111011000100001000100010011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100001110111011101111000100001110111011001100101010101000100010001000100010001000100001100110011001100110010001000100010001000110011010001000011001000110100010001010100010000110010001000100010001000100010001000100010001000100010001000100011001100110011001101000101011001111000011110000111011101100101011001110111011101010100010001000101011001111000100010011001100110011001100110011001100110011001100110000111010101000100010001010101010101010101010101010110011101110111100010001000100001110100001101000100001100110011001100110011001100110011001100110011001100110100010001000101010101010101010101000101010001010110011101100110011101110111011101111000100110011001100110011001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100110011001100010001000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110101000100010001000100110111100001110111011101111000100010001000100001110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011101110111010000100001000100100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000011101110110011001010100010001000100010001000100001100110100001100110011001100110011001100110011001000100010001000100010001000100010001000100011001101000100001100110010001000100010001000100010001000100010001000100010001000100011001100110011001100110100010101010111011101111000100001110101011001110111011101010100010001000101011110001000100110011001100110011001100110011001100110011001100001110110010101000100010001010101010101010110010101101000011101111000100010011000100001000011010001000100001100110011001100110011001100110011001100110011001100110011010001000101010101010101010101010101010001010110011101100110011101111000011101110111100010011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000011101110111011101110111011101110111011101110111011101111000100010001000011101110111011101110101001000010001000100100110100010001000100010001000100010001000100010000111100010001000011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111100001110110001100100001000100100101011110000111100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000100010001000100010001000100001110110010101000100010001000101010101000100001100110011001101000100010001000100001100110100010001000011001100100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110100010001010101010101101000100001110110011101110111011101000100010001010110011110001000100110011001100110011001100110011001100110011001100001100101010101010100010101010110011001100110011001111000100010001000100110010111010101000100010101000100001100110011001100110011001100110011001101000011001100110011010001000100010101010101010101010100010101010110011001100110011001111000100010001000011110001001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010000100100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000011101110111011110000101001000010001000100100110100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101111000100010001000100001110110001000010001000100100101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000100010000111011101010100010001000101010101010101010101000100010001000100010001010101010101010101010001010101010101010100001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011010001000100010001000011010001000101010101010100010101101000100010000111011101111000011101000100010101010110011110001001100110011001100110011001100110011001100110011001011101100101010101010101010101010110011110000110011110001001100110011001100001110110010001010101010101010011001100110011001100110011001100110011001101000011001100110011001101000100010101010101010101010101010101010110011001110110011001111000100010001000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100001111000011101110111011101110111100010000111011101110111011110000110001000010001000100100110100001111000011101111000011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011110001000100010001000100010001000100001110101001000010001000100110110011101111000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110100010001000100010001000100010000111010101010101010101010101010101010101010101010101010101010101011001100110011001100101010001100110011001100101010001000100010001000011001000100010001000100010001100110011001000100010001000100010001000100010001000100010001000110011001100110011010001010101010101100110011101110110011001101000100010000111011110001000011001000100010101010111100010011001100110011001100110011001100110011001100110011000011001100110011001010101011001100111100010010110100010011001100101110101010001000101010101010110011001000011001100110011001100110011001100110011010001000011001100110011010001000100010001010110011001010101010101010101011001110110010101101000100110011000100010001000100010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010001000100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001110111011101110111011110000111100001110111011101110110001000010001000100100101011101110111011101110111011101110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100010000111011101110100001000010001000100110110011101111000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100001110110011001100101010101100110011001100110011001100110011001100111011101110111011101110110010101100111011101100110010101010101010000110010001000100010001000110011010000110011001000100010001000100010001000100010001000100011001100110011001100110011001100110011001101000101011001110111011101111000100101110101011110001000010101000100010101100111100010011001100110011001100110011001100110011001100110011000011001100111011001100110011001111000100110011000100010011000011001010101010101010101010101010110011001000011001100110011001100110011001100110011010101000011001100110011001101000100010001000101011001100101010101010101011001110110011001101000100110011001100010001000100010001001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001110111011101110111011110001000011101111000011101110111001000010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100001110111011101110011000100010001001001010111011101111000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110110011001110111011101100110011001100101001100100010001000100011001101000100010000110010001000100010001000100010001000100010001000100011010001000100001100110011001100100011001100110011010001100111011001111000100001100101011010001000010101000101010101101000100110011001100110011001100110011001100110011001100110011000011101110111011101110111011110001001101010101001100010000101010101010101010101010101010101100111011001000100010000110011001100110011001100110011010101000100001100110011001101000100010001000101011001100110010101010101011001110111011001101000100110011001100110001000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001111000011101110111011101110111100010001000011101110111011101110111001100010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100001110111011101100011000100010001001001010111011101111000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100111100010001000100010001000011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100110010101000011001000100010001000110011010001000100010000110010001000100010001000100010001000100010001000100011001101000101010101000011001100100010001000110011001101000101010101100111011001000101011110001000010101000101011001111000100110011001100110011001100110101010100110011001100110101000011110001000100010001000100110011010101010101010100001010101010101010101010001000101011001100111010101000100010000110011001100110011001100110011010001000100001100110011001101000100010001000100010101100110011001010110011001100111011101100111100110011001100110001000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000011101110111011101111000100010000111011101111000011101110111010000010001000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100001110111011101010010000100100010001101010111011110001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101101000100010001000100010000111010101100110011101110111011101110111011101110111100001111000011101110111011101111000100001110110011101110111011101100110010000100010001000100011001100110100010001010100001100100010001000100010001000100010001000100010001000100010001100110100010101010100001100110011001000100010001000110011001101000100010001000100011110000111010001010101011001111001100110011001100110011001100110101010100110011001100110101001100010011001100110011001100110101010101010101001011001010101010101010100010101010110011101110110010001000101010000110011001100110011001100110011001101000100001100110011001100110100010001000100010001010110011001100110011001110111011101110111100110101001100110001000100010001001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101111000100001110111011101111000011101110111010000010001000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010000111011101110111011101000010000100100010010001100111011110001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101101000100010001000100010000110010101100111011101110111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101010011001100100010001000110011001101000100010101010011001000100010001000100010001000100010001000100010001100100010001000110011010001010101010000110011001000100010001000100011001100110011001100110100010101110110010001010101011010001001101010011001100110011010100110011001100110011001100110101001100110101010100110101010101010101010101010100111010101010100010101010101010101100111100010000101010001010101010000110011001100110011001100110011010001000100001100110011001100110100010001000100010001000101011101110110011001111000011101110111100110011001100001111000100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000100010000111011110000111011101110111010000010001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011110001000011101110111011101110111011100110001000100010010010101110111011110001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000100010001000100001110110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010000111011101110111010100110011001000100010001101000100010001000100010000110010001000100010001000100010001000100010001000100010001000100010001000100011001101000100010001000011001100100010001000100010001000110011001100110100010101110101010001010110011010011001100110011001101010011001100110011001100110011001101010101010100110101010101010101010101010101010101010010110010101010101010101010101011001111000100110000100010001100101010000110011001100110011001100110011010001000100001101000100001100110100010001000100010001000100011001110111011001111000011101110111100010011001011101100111100110011001100110001000100110101010101010101010101010101010101010101010101010101010101110111011101110111010101010101010101010101010101010111010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110101001100110011001100110011001100110011001100001000010000100100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110000111011101111000011101110111011101111000010100100001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011000100001000100100011010101110111011101111000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000100010001000100001110111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110101001100100010001000100011001101000100010000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011010001000100001100110010001000100010001000110011001100110100010001100101010001010110011110011001100110011001100010001001100110011001101010101010101010101010101010101010101010101010101010101010101001110101010101010101010101010110011110001001100101100100010101010100010000110011001100110011001100110011010001000100010001000100010000110100010001010101010101000100010101100111011001111000011101110110011110011000010101010111011101110110011001111000100110101010101010101011101110111011101110111011101110111011101110111011101110111011101010111010101010111010101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011010100110011001100110011001100000110001000100101000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110000111011110000111011101110111011101110111011101111000011000100001000100010001010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111010000100001000100100011011010000111011101111000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001000011001000100010001000110011001100110100010001000100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001101000100001100110011001000100010001000100011001100110100010001000100010101010101011110011001100110011000011101111001100110101010101010101010101010101010101010101010101010101010101010101011100101100101010101010101010101100111100010101010100001000100010001000011010001000100001100110011001100110100010001000100010001000100010000110100010001010110010101010100010101010110011101100111100001110110011110010111010101010110010101010101011001111001100110101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001101010101010101010011001100110011001100000110010000100101000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100001110111011101111000011101110111011101110111011000100001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111001100010001000100100011011010000111100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100100001100110011001000100010001100110011001100110100010001000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010000110011001100100010001000100010001100110100010001000100010101010101100010001001100001110111100010011001101010101010101010101010101010101010101010101010101010101010101110101010011101010101010101010101011001111000100110101010011101000100010001000100010001000011001100110011001101000100010001000100010001000100010001000011010001000101010101010101010101010101011001110111100001110110011010000111010101010101010101010110011110001001101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010100000110010000100111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101111000100010001000100001110111011101110111011000100001000100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110110001000010001000100100100011110001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101000011001100110011001100110011001100110011001101000100001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001000011001100110010001000100010001100110011010001000100010101010101011010001000011001111001100110011010101010101010101010101010101010101010101110111011101110111011101110111000010101010101010101010101011001111000101010111001010101000100010001000100010001000011001100110011001101000100010001000100010001000100010101000100010001000101010101100101010101010101011001110111100001110101010101110101010001010100010101010110011110001001101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000110010000100111000101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010000111100001110111011101111000011100110001000100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110100001000010010001000100101100001111000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110101001100110100001100110011001000100011001000100011001100110011001100110011001000100010001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001100110011001100110011001000100010001000110011001100110101010101000100011001100110011110011001100110011001101010101010101010101010101010101011101110111011101111001100110010110111010101010101010001010101011010001001101010111000010001000100010001000100010001000011001100110011001101000100010001000100010001000101010101010100010001010101010101010101010101010101010101100111100010000101010001100101010001000100010001010110011110001010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000110010000100111000101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100001110111011101110111011101111000011101000001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110011000100010001001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010100001101000101010000110011001000110011001000110011001100110011001100110011001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100100010001000110011001101000100010001000100010001010101011001111000100110011001101010101010101010101010101110111011101110111011101111001011101110000101010101010101010101010110011110011010101010100110010001000100010001000100010101000100001100110011010001000100010001010101010001010101011001100100010101100101010101010110011001100101010101010111100001110110010001000100010001000100010101100111100010011010101010101010100110011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000110010000100111000101010011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101000001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101010010000100010001001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000100010001000100010001000100010001000100010001000100010001000100001110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000100010001010100010000110011001100110011001100110011010001000100010000110010001000100010001000100010001000100010001100110011001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110010001000110011001101000100010001000100010001000101010101100111100010011001100110101010100110011001100110011010101010101010101110111011101001100101010101000100010101010111100110101010101110100101010001010101010101010101010101000100010000110100010001000100010001100110010101010110011101110101010101110111011001010110011101100110011001010110011110000110010001000100010001000101011001111000100010011001100001110111100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000100010000100111000101010101010101010101010100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100010011001100110001000100010001000100010001000100010001000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111100001010010000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101000010000100010001001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000100010101100101010000110011001100110011001100110011010001000100010000110010001000100010001000100010001000100011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001101000100010001000100010001000101010101100110011101111000100010001000011110001000100110011001100110101010101010111011100101100101010101000100010101100111100110111011110010100101010101100101010101010101010101000100010001000100010001010100010101110110011001100111100010000110010110001001100001110110011001100110011001100110011110000110010001000100001101000110011110001000100010001000011101111000101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110010111100101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010100000100010000100111001101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010011000100110001000100010001000100110011001100110001001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011000110010000100010001001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010001000100010001000100010001000100010001000100001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010001000101011001100110010000110011001100110011001100110100010001000100010000110010001000100010001000100010001100100011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001101000100010001000100010101010101011001110111011101111000100010001001101010101011101110111011101110111011100101010110011001000101010101101000101010111100110010000101011001100110010101010101010101010100010001000100010101010100011010000111011101111000100110010111010110011011101010011000011101100110011001100111011101110101010000110011010001010111011101110111011001100111100010101010101010111011101110111011101110111011101110111011101110111011101111001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110001001100110011001100110011000100010001000100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011000100001000100010010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010001000100010001000100010001000100010001000100001100111100110001000100010001000100010001000100010011001100110011001100010011001100110011001100110011000100001110101010001010101011001100101010000110011001100110011001100110100010101010101010000110011001000100010001000100010001100110011001100110011001000100011001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110100010001000100010101010110011101110111011101110111100010011001100110011010101010111011110010111011100101010110011001010110011001111001101111001100110001110101011101100110011001100110010101010100010001000100010001000101011110001000100010001001101010101000011010011011101010101010100110000110011001100110011001100100010000110011010001100111011001100110011001100110100010101010100110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011000100010001000100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011000100010001000100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111010000100001000100010010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000100001101000100110001000100010001000100010001001100110011001100110011001100010011001100110011001100110011001100001100100010101010101011001010101001100110011001100110011001100110101011001100101010000110011001100110010001000100010001100110100010000110011001000110100001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001000100011001100110011001101000100011001111000100001110111011110001000100010011010101010101011101110111011101110111011100001010111011001010111011101111010101111001100101101010110100101110111011001100110010101000100010001000100010001010101011101111001100110011010101010101001011010011011101010101001100010000111011101100101010101010100001100110011010101100110010101010101011001101000100110111011101010111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100110011001100110011001100010011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011000100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111001100010001000100010010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000100001101000100110011000100010011001100110011001100110011001100110011001100110011001100110011001100010011001011101010101010101010110011001100100001100110011001100110100001100110110011101110101010000110011001100110011001000100010001101000100010001000011001001000101001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110010001100110011001101000110011010001001100101110110011110001000100010011001101010111011110011001100110011001011100001010111100001101000100110001011110011001101101001011000100110000111011101110110010101010100010001000100010001010110100001111001101010101010101010111001011010001010101010111010100110000111100001110110011001000100001100110100010101100101010101010101011001101000100110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100000100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110110001000010001000100100011010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001001011101101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011001000100010001010110011101100101001100110011001100110100010001000110100001110101010000110011001100110011001100100010010001010101010101000011001101100101001100110011001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001101010110011101110111011001110110011001100111100010001000100110101011110011001100110011001100100001011000100001111010101010101100110111001101100101011001101010011000100001110111011001010100010001000100010001010111100001101010101110111011101110101000011001111001100110011001100110011000011101110110011001010011001100110100010101010110011001100110011001110111011110011010101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100110011001100101110111011101110111100110011001011101110111011101110111011101110111011101111001011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100000100010001001000100101011101110111011101110111011101110111011101110111100010000111011101110111011101110111011101110111100001110111011101110111,
	2400'b011101110111011101110101001000010001001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001011101111000100010001000100010001000100010001000100010001000100010011000011001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111010101000100010101010110011101110101001100110011001100110011010001000110100101110101010001000011001100110011001100100010010101110111010100110011001101110110010000110011001100100010001000100010001000100010001000100010001000100011001100110011001100110011001101000100010000110100010001000101010101100110010101010101011001110111100010001001100110101011101111001100110011001100100101101001101010001011101110111101110111011101100001101011100110001001100110001000011001010101010001000100010001011000100101101001110011011011101110101000011101110111011101100110011001100110010101010100010001000100001100110100010001010110011001110111100010001001100110001000100110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111001100110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101000100010010001000010100011101110111011101110111100010001000100010000111011101110111011101110111011101111000100010000111011101110111011101110111,
	2400'b011101110111011101110011000100010001001000100100011110001000100010001000100010001001100010011000100010001000100010001000100010001000100010001001011101101000100010001000100010001001100010001000100010001000100110011000010110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000110010101000100010001000110011101100100001100110011001100110100010001011000100101100101010001000011001100110011001100110011010001110111010000110011010001110111010100110011001100100010001000100010001000100010001000100010001000100010001100110011001100110011001100110100010001000100010001000100010001010101010001010101011001110111100010011001101010111011101111001100110011001100100101101001101010011100110011001101110111011100011010001011101010011010101010011001011001010100010001000100010001011000100001011001110011001010100110101001011101100110011001100101010101010101010101010100010001000011001100110011010001010110011101110111100110011010101010101010100010001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011100000100010000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100110001000100110011001100110011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000010001001000010011011101110111011110001000100010001000100010001000100001110111011101110111011110001000100010001000011101110111011101110111,
	2400'b011101110110011101100010000100010001001000110101100010001000100010001001100110011001100110011001100110011000100010011001100110011001100110001001100001101000100110011000100010001000100010001001100110011001100110011000010110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100101010001000100010101010110011001010011001100110011001101000100010001011000100101100101010001000100001100110011001100110011001101000100001100110011010010001001011000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011010000110011001100110100010001000100010101010101010101100110011110001001101010111011101111001100110011001100101001111010101110101101110111011101110111011100011010011100101110111011101110111010011101100101010001000100010101101001011101011000110011001011100001110111011001100110011001100110011101110110010101000100010001000100010001000100010001000110011001111000100010011010101110111011101110011001110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011001100110011001100110011001100110011001100110011001100110011001100110111001101110111011100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011100000100010000100111001101110101011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000010001000100010011011101110111100001111000100010001000100010001000100001110111011101110111011110001000100010001000100001110111011101110111,
	2400'b011101110110011101010010001000010010001000110110100110001001100010011001100110011001100110011001100110001000100010011001100110011001100110011001100001101000100110011001100110011001100110011001100110011001100110011000010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001010100010001010101010101010110010000110011001100110011010001010101010101101001100101110101010001000100010000110011001100110011001100110011001100110011010001111000011001000011001100110010001000100010001000100010001000100010001000100010001000100010001100100011001000110011001100110011001100110100010001000100010001000100010001010101010101100111100010011010101110111011101111001100101001111010101110101101110111011101110111011011010110101100101111001100110010111011100101100101010001000100010001111010011101011001101010111100101110000111011101101000100010001000100001100101010001000100010001000100010000110011010001000100010001010110100010001010101110111100101110111010101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011100000100010000100111001101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100010001000100010010011001111000100001111000100010001000100010001000100001110111011101110111011110001000100010001000011101110111011101110111,
	2400'b011101110111011000110010001000010010001101000111100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001101000100110011001100110011001100110011001100110011001100110010111011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011001000101010101100110010101010101010000110011001100110011010001100110011001111010101001110101010101000100010001000100010000110011001101000100011001100100010001111000011101000011001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010101000100001100110011001100110100010001000100010001000100010001010101010101100110011110001010101111001100101010001010110010111101110111011101110111011001010110111100110011001100110011001011100101100101010001000100010110001010011001101001100110011010100110000111011101111000100010001001011101000100010001000100010001000100010000110011010001000100010001000101011001111000101010111100101110111100101111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111100101110111011101110111011101110111011100000100010000100111001101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100010001000100010010011001111000100010001000100010001000100010000111011101110111011101110111011110000111011110001000011101110111011101110111,
	2400'b011101110111011000110010001000100010001101011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101101000100110011001100110011001100110011001100110011001100110010110011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011001000110011110000110010001000011001100110011001101000100010101110111100010011011101010000101010001000100010101010101010000110011010101110110100001010100011001111000011000110011001100100010001000100010001000100010001000100010001000100010001000100011001100110011001100110100010001000100001100110011001100110011001100110100010001000100010001000100010101000101010101100111101010111011101010001011110010111101110111011101110111011000011111001100110011001100110010111011100101110101010101010100010110011010011001101001100110011001100010001000011101110111011110010111010101000100010001000100010001000100001100110011010001000100010001010101010101100110011110001010101111001100110010111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111100101110111011101110111011100000100010000100111001101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000010001000100010001010101110111100010001000100010001000100010001000100010001000011101110111011110001000100010001000011101110111011101110111,
	2400'b011101110111010000100010001000100010010001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100110011001100110011001100110011001100110011001100110010110011110011001100110011001100110011001100110011001100110101010101010101010101010101010101010011000011001101000100110000101010101000011001100110100010001000100011001111000100010101011101010000110010101010101010101100111011001000011011010000110011101000101010101100101010000110011001100110011001100110011001000100010001000100010001000100010001000100011001100110011001100110011001101000100010001000100010000110100010001000100010001000100010001000100010001010101011001100111100110111011101010011011110011001101110111011101110111010110100011001100110011001100110010111011101001110101010101010100011010101010010101101001100110011001101010101001011101101000100101110100010001000100010001000011001100110011001100110011010001000100010001000101010101010110011110001000101011001101110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011011100110011011101110011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100100000100010000100111001101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100001000100010001010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011101110110010000100010001000100011010110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100110011001100110011001100110011001100110011001100110000101100010101001100110011001100110011010101010101010101010101010101010101010101010101010101010101000011110001001100001100101010101000011001101000100010101010110011010001001100110101011101110010111011001110111011110001000011001000011011101100101010101000101010001000100010101010100010000110011001100110011001000100010001000100010001000100010001000100010001000100011001100110011001100110011010001000100010001000100010001000100010001000100010001000101010101010110011001100111100110111011101010101011110011001101111011101101110111000110101011001100110011001100110011001100101001110110011001010101011110111010010101111010100110011010101010101001011110001001011001010100010001000100001100110011010000110011001100110100010001000100010001000101011001110111011110001000100010011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100100000100010000100111001101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000010100100001000100010001001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011101110110001100100010001000100011011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000110100110011001100110011001100110011001100110011001100110000101100110101001100110011010101010101010101010101010101010101010101010101010101010101010101010101000100010001000011001010101010101000011010001000100011001111000100010001010101010111011101110101000100010001000100010001000010100110011011001000100001100110011010001000101011001100101010001000100001100110011001100100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110100010001000100010101010101010101010110011001100110011110000111100110111011101010101011110011011110111011101101111010110110101111001100110011001100110011001100101101110111011101010101100111001010010110001010101010101011101110111001100110100110010101000100010001000100010001000100001100110100010001000100010001000100010001000100010101111000100010001000100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010000100111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000011000100001001000010001001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011101110100001000100010001000100011011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000110100110011001100110011001100110011001100110011001100101110110100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100001110111011101100101010101000100010001000101011110001001100110011010101110111011101110101000100110001001100110000111010000100011010000110011001100110011010001010101010101010100010001000011010000110011001100110011001000100010001000100011001000100010001000100011001100110011001101000100010001010101010001010100010001000100010001010110100010001000100110011001100110111001100110101011101010111011110011011110111011101110110110010110110011001100110111011101110111011100101010000111011001010101101011011010010110001011101110111011110010111011101001110101010001000100010001000100010001000100010001000100010001000100010101010100010101010101010101010111101010101010100110101001100010101100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110111011100110011001100110011001100110111011101110111011101110111011101110111011100110111011101110011001100110011001100110011001100110011001100110011001100110011001100100000100010000100111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000011000100001000100100001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011101100011001000100010001000100011011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110100010011001100110011001100110011001100110011001100101100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010111011001111001100001010101010101000100010001000110011110101011101110111011101110111011101110111010101010101010100101110100001100100011001100110011001101000100010001000100001100110011001100110011001100110011001100110011001100110010001000100010001000100010001000100010001100110011010001000101011001110111011110001000011101110111011001100110100010101011101111001100110011001100101110011001101111001100110111011110111011101110110101111000110111001100110111011101110111011100101110001000011001010110101111011001010110011011110011001100110011001100100001100101010001000100010001000100010001000100010001000100010001000100010101010101010101100101010101010110100110111011101110101010100110011011110111011101110111011101110111011110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100100000100010000100111001110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000011100100001000100010001001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011101010001001000010001001000110100011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110100010011001100110011001100110011001100110011001100101100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010110011110011001011001010101010101010100010001000110100010101011101110111011101111001011101110111011101110111010100001000011001000100011001100100011001101000011001100110011001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000100010001100110011001100110100010001010110011110001001100110011001100110011000011001101001101111001100110111001100110010111010101010111100110111101110111011101110110001101010110111001100110111011101110111011100101010011001011001011000110111011001010110101100110011011101110011001000011001010101010001000100010001000100010101100101010001000100010001000100010001100110010101100110010101010110011110111100110011001010101010101010110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011110110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100100000100010000100111001110010111100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011010100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000011100110001000100100001001001010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011000110001000100010010001101000110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011110011001100110011001100110011001100110011001100101011000101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110011000100110101001011001010101011001010101010001000110100110101011101110111100110011001011101111001011101110101000010000110010001000100011001100100011001100110011001000100010001000100010001000100010001000100010001100100010001000100010001000100010001000100010001000100011001100110011001100110011001101000100010101100111011110000111011110001000100001100110011110011011110011001100110111011100101110111100110111101110111011101110101001101100110111011101110111011101110111011101101110111001011001011010110111011000011011001101110111011101110110100111011001010101010001010101010001000101011001100100010001000100010001000100010001100111010101100111011001100110011010011100110111011100101110101011101111001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110110111011110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110110111101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100100000100010001000111001110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100001000001000100010001000101000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b011000100001000100010010001101011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011010011001100110011001100110011001100110011001100001011001101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110101010101010100111011001010111011001100110010101100111100110111011101110111100110011001011110011001011101110000101001100100010001000100011001100100011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001000011001100110011010001000100010101010101010101010101011001100101010101010111100110111100110011011101110111001100110111101110111011101110100001111101110111011101110111011101110111011101110111001001010101101100111011010111011111011101110111011101110010011000011001010100010001100101010001010110011001010100010001000101010101000100010001101001011101010111011101110111011001111010110111011101110111001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100100000100010001000111001110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100001000001000100010001000100110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b010100100010000100100010001101101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011010011001100110011001100110011001100110011001011101011001101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111010101010010110010101111000011101110111011110000111100110111100110011001100110011001011110011001011100101100101001100100010001000100011001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010001000100010001000100010001010110011001010101010101000100010101010110011010001010110011011101110111011101110111101110111011101101011010011101110111011101110111011110111011011110110111011000010101111101111011010111100011011101110111101101101110101000011001010101011001100101010101100110010101000100010001000101010101010101010001011001101001110111100010000111011110001001101111011101110111011101110111001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111101111111111111111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100100100100010001000111001110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100001010001000100100010000100100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100010001000100100010010010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010110011001100110011001100110011001100110011001011001101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101001110110011010011010100010001000100010101001101010111100110011001100110011001100110010111010100101110100001000100010001000100011001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001100110011001100110100010001000100010001000100010101100110011110000111011001010100010101010101011001111001101011001101110111101110111011101110111011101100011010111101110111101110111011101110111011101110111011000111010110101110111011010110100111011110111011101110110010101000011001010110011101100101011001100101010001000100010001010110011001010101010101010111101010000111100110011000100010001001100111001110111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100100100100010001000111001110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100001010001000100010001000100100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001000100100011010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010110001001100110011001100110011001100110011001010101111010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110101001100001111000100110101010100010001001101010111011101010111100110011001100110011001100110010111010100001000011001000100010001000110011001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001000100010001000101010101100110011001111000100010000101010001010101010101101000100010111100110111011110111011101110111011101001011011001101110111101110111011101110111011101110111011000110011011001110111011000110101111101110111011101110110110111000011101101000011101100110011001010101010001010101010101100111011001100110010101000101100010011000100110101010100110011010101010101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100100100100010001000111001110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011010101010011001100110011001100110011001100110011001100110011001100110011001100010001000100101100010000100010001000100100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001001000110100011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010101111001100110011001100110011001100110011001010110001010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110101000100010001010101110111011100110001010101111001100101110111100110011001100110011001100110010111000010000110010001000100010001000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110100010001000100010001010111100001100111100010100111010101010110011001100111011110001001101111011110111011101110111011100111100011011101110111101110111011101110111011101110111010110110100111011110111010110110110011101110111011101110110110111001100010001001100001110110010101010101010101010101010101100111011101110110010101010100011110101001100111001100101110101011101110011011111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111101101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110011001100110010111011100000100010001000111001110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110001000100101110010000100010010000100010100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001001001000101011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101111001100110011001100110011001100110011000010110011010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111010011110101011101111001011101010011011101111001100110011001100110011001100110011001100101101110100010000110010001000100010001000110011001100110010001000100010001000100010001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001101000100010001000101011110001000100110011001100001100111100010001000100010001000100010101100110111101110111011000101101011011101110111101110111011101110111011101110111010010110101111101110111010100111110111101110111011101110110111001010100010101010100110000110010101010101010101010101010110001000011101110111011001010101011010011011100111001110110111001011110010111010110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111001100101110111011101010101010011100100010001000111000101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100101110010000100010010001000010011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001001001000101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001010101101001100110011001100110011001100110010111010110101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011110011001011101010111100110011001100101010011011110011001100110011001100110011001100110011001011011101000101001100100010001000100010001000110011010000110010001000100010001000110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110100010001000100010101101000101010011000101010000111100110011010101010101001100010011001101111011110111010010101110011011101110111011110111011101110111011101110111001110111110111101110111010011000111011101110111011101110111011011011100110111011101010010110010101010101011001100110011010011000011110000111011001100101010110001100101110111110110111011100110111001001101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111001100101110111010101010101010101010101010011100100010001000111000101010101010101010101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101011101110101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110000011000100010010001000010011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010010001101000110100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011000011101111001011001101001100110011001100110011001100110010111011010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011110011001100101111001100110011001100101010101100110011001100110011001100110011001100110011001000010101010100001100100010001000100010001000110011001100110010001000100010001101000101010000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001000100010001000101011110011001101110101001101010101011110011001011101010101010101010101101111001100111110111011101110111011110111011101110111011101110110101111001111011101110111010001001111011101110111011101110111011011100101010111100101110010101010101010101011001100110011110011001011110001000011101100101010101111100110010111101111011011101110111001001100010111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111001100101110111010101010101010101010101010101010101010011100100010001000111000101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010010100000100010001000100010010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100100010001101000111100010001001100110011001100110011001100110011001100110011001100110011001010101000101011110001001100110011001100101100100001100110110011101111001100110011001100110011001100110010110011110101010101010101010101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100101110111100110011001100110011001100110011001100110010010110011001000011001100100010001000100010001000110011001100110010001000100011001101000100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001000100010001000100010001101000101010111010101011001100110011011100110011001011101110101011101101011010110111011101110111101110111011101110111011101110101101101011111011101110111001111010111011101110111011101110111011101100101010101011101101110101010101100110011001101000011110101001100010011001100001110110010101101100111011011101111011011101111011011010100110011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001011101110111010101010111011101110111011101110101010101010101010011100100010001000101000101110101010101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110101011101110111011101110111011101110111011101110111011101110111011101110111010101110111011101110111011101110111011101010101010101010100110000100010010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100100011001101010110010101011000100110000111011010011001100110011001100110011001100110010111010000110100010001000101011110011010100101010011010001000100010001011001100110011001100110011001100110010101100010101011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100101110111100110011001100110011001100110011001100110010010111010001000011001100100011001000100010001000110100001100110010001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110100010001000100010001000100010001010101011110101011101011001101110111011101110111001100110010111011100001011011110111011101110111101110111011101110111011101110100101101101111011101110110101111100111011101110111011101110111011101101101110011010100001111000011001111000011101101001100010011000100110011001100001110110011001101011111011101101111011011110111011101011100110001100111111101111111111111111111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001011101110111011101110111011101110111011101110111011101110111010101010101010011100100010001000101000101110101011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010100110011001100110010111001000010001000100100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011001101010100001100110101010101010100010001101001100110000111011101111000100110000100001101000100001100110011001101101000100001110100001100110011001101000111100001110111100010011001011101010100011010011011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110000110010101000011001100110010001000100010001101000011001100110011001100110011001100100010001000100010001000100010001000100010001000100011001100100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001000100010001010101010101010101010101101000101011001101110111011101110111011101110011001011010101101011101111001101110111011110111011101110111011101110011110001110111011101111110001111101111011101110111011101110111011101101110010101001100010001001011101111000011010011010011110011001100110101001100110000110011001101010111011101110111011101110111111101100100110011101111111111111111111101111111111101110111111111111111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001011101110111011101110111011101110111011101110111011101110111011101110111011101010101011011100100010001000101000101110101011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010111011101110111011101110111010101010101010101010101010101010101010101010101010100110011001100110011001100010001000100010000111001100010001000100100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001101000011001100110011001100110011001101001000100101100100010001000101011101110011001100110011001100110011001100110011010101100100001100110011001100110100010001000011010001100110010000110011011010101011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011011100110011001100110011001100100101110101010101000100010000110011001000100010001101000011010000110011001100110011001000100010001000100010001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011010001000101010101010101010101010110010101010101011110011100110111011101110111011101110111011011010010001011101110111011110011001101110111101110111011101101011010101110111011101111101110001110111011101110111111111110111011101110110110111001100110011001011110000110011111001101100010101011101010011010101010010111011001101010111011101110111011101110111111101100101010011101111111111111111111111111111111111111111111111111111011101111111111111111111111111111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111011111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011011100100010001000101000101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010000111001100010010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010010001000010001000110010001100110011001101000101011001010011001000100011010101000011001000110010001000100011001100100011001101000011001100110011001100110011001100110011001101000100010000110100101010111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011011101110111011101110011011101110011011100110011011100110011001011100001100100010101010100001100110011001000100011001101000100010000110011001100100010001000100010001000100010001000100010001000100010001101000011001100100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001101000101010101010101010101010110011001010110010101101001110011011101110111011110111011101010010110101011101110111011101110111011110011001101111011101011010111001110111011101111100110011110111011111111111111111110111011101110110110111001101010111010011101110110110011101101100010111101110010111100101110101000011001101010111011101110111011101110111111101101101110101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100000100010001000101000101110101011101110111011101110111011101110111011101110111010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000010000010010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011010000110010001000100010001100110011001100110101010000110011001000100010001100110010001000100010001000110011001100100010001100110011001100110011001100110011001100110011001100110100010000110110101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110011001010011001010101011001000011001100110011001100110011010001000100001100110011001000100010001000110011001000100010001000100010001000100010001101000011001000100010001000100010001000100010001000100010001000100010001100110100010000110011001100110011001101000101011001100110011001100110011001100110011001100110100111011110111011101110111011101000011011001101110011001011101110111011101110111011110011011000011011011110111011101110100010101110111011101110111111111110111011101110110111001011110011011011011101101001111011101101100011011110111011011100110010111001011101111010111011111110111011101110111111101110111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100000100010001000100111101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101011101110111011101110111011101110111011101110111011101110111010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000010100100001000100100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011010000110010001000100010001000100010001000100011010000110010001000100010001000100010001000100010001100110010001000100010001100110011001100110011001100110011001100110011001100110100001100110111101110111011101010111011101110111011110010111011101111001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111001000011001100110010101000011001100110011001100110011010000110011001100110011001100110011001100110010001000100010001000100010001000100011010001000011001000100010001000100010001000100010001000100010001000100010001000110100010001000100010001000100010001000100010101110111011101110110011101100110011001100110011110111110111011101110111011010110100011011101110111011101110011001100101110111011101110110110100011011101110111101101011110111111111111111111111111111110111011101110111011011101110111101011011101111101111011111011100111101110111011101101110011001010100010001010111011111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100000100010001000100111101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000011000100001000100100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011010000100010001000100010001000100010001000100011001100110011001000100010001000110011001000100010001100110011001000100010001100110011001100110011001100110011001100110011001100110011001100110111100110100111011001110110011001111001101110111011110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111001000011001110110010101000100001100110011001100110011001100110011001100110011001100110011001100110010001000110011001100100010001000110100010001000011001000100010001000100010001000100010001000100011001000100010001000110100010001000100010001000100010001000100010001101000100010001000100010000111011101100111011110001100111011101110111011000100101011011101110111011101110111011101110010111011101110100100100111011101110111011011011111001111111011101110111011101110111011101110111011101110111011101011011010101110111011101010101111101110111011101101110111011011100110011010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111011111111111111111111111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100000110010001000100111101110101011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000011000100001001000100010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011001100100010001000100010001000100010001000100011001100110011001000100010001000110011001000100010001100110011001000100010001100110011001100110011001100110011001100110011001100110011001100110110100001010101011001100011001101000101101111001100110010111011101111001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110110111000011101110110010101010100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100100010001101000101010101000011001100110011001000100010001000100010001000100011001000100010001000110011010001000100010101000100010101000100010001000110100110101010101010011001100010000111011101111001110111101110111010010101110011011101110111011101110111011101110111011100110010010100101111011101110111011010011111011110111011101110111011101110111011101110111011101110111011101001011111001111111011101000110111101110111011101110110111011100101110111011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111110111011111110111011111111111011101111111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100110010001000100111101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000011100110001000100100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011001100100010001000100010001000100010001000100010001100110011001100100010001001000011001000100011001100110011001000100010001100110011001100110011001100110011001100110011001100110011001101000111011001010110010101000011001100110101100110011001100001100110011110101011110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110110111000100001110101010001010101010101010101001100110011001100110100010001000100001100110011001100110011010001000011001100110010001101010110011001000011001100110011001000100010001000110010001000100011001100100010001000110011010001000101010001010101010101010101010001000100011110111011101110101010101010101001100010001000101011101110111001110110110111011101111011101101110111011101111011011101111010000101110011011101110111011001011111011101110111011110111011101110111011101110111011101110111011101000100111101110111111001000111011101110111111101110111011101101110011001100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011111110111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100110010001000100110101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110011001100010001000100010001000100001000001000100100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011001100100010001000100010001000100010001000100010001000110100001100100010001000110011001000100011001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110100010001000100001100110011001100110011010001000100001100110011010001011001110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110110101001100101110110010101110111011001100100001100110010001100110101010101000100001100110011001100110100010101010011001100110011010101110111010100110011001100110011001100100010001100110010001000100011001100100010001000110011001101000100010001010101010101010101010001010100010110001011110011001011110011001011100110011000100011001110110001011000111011101110111011101110111011101110111011011110110101100111110111011101110111010111100111011101110111011110111011101110111011101110111011101110111111000111110011111110111110101001111011101110111011101110111011101110111011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111110111011111110111011111110111011101110111011101110111011101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100110010001000100110101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100001010010001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011001000100010001000100010001000100010001000100010001000110100010000110010001000110011001000100010001100100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000110011001100110011001101011001110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110010111011100110000111100010011000100001010011001100110011001101000110011001010100001100110011001101000110011001010011001100110101011110000110010000110011001100110011001100100010001100110010001000100011001100110010001000110011001101000100010001000101011001100110010101010101010001011000101111001100110111001100101110011011100110011101100101001010111011101110111011101110111011101110111011101110110101011001111011101101110111010110101011011101111011101110111011101110111011111111111111101111111110101000110111111110111010001011111111101110111011101110111011101110111011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111110111011101110111011101110111111101110111011101110111011101110111011101110111011101111111011101110111011011101110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100110010001000100110101010111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100001100010001000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100011001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001101010110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110011001011101010101001101010111011011100110011001100110011001101010110011001010100001100110011001101010111011101000011001101000111100001110100010001000011001100110011001100100011010001000010001000100011001100110010001000110011010001000100010001000101011001100110011001100101010101010101100010111100110011011101110010101010101110011011011001011100111011101110111011101110111011101110111011101110101101011011111011101110111011000110101111101110111011101110111011101110111011111110111111111111111010001010111111111110110001111101111111101111111011101111111111101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111101110111011101110111111111111111011101110111011101110111011101110111011101110111011101101110111001100110011001011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100110010001000100101101010111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001100010001000100010001000100001110011001000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100001000100100010001000100010001000100010001000100010001000100010001000110011001000100010001000100010001000110100010000110011001100100011001100110011001100110011001000110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011010110001000100001110111100111001100110011001101110111011101110111011101110111011101110111011101110111011101110111001011101110111011110011001010010100110011001100110011001101000110010101000011001100110011010101111000011001000011010001101000011101010100010001000011001100110011001100110011010001000010001000110100001100110011001100110011010001000100010001000110011001110110011001100101010101010101010110001011110011001101110010111010101010010111010001101101111011101110111011101110111011101110111011101110100101011101111011101110111010110110110111101110111011101110111111111111111011111111111111111111110101111100111111101110101010011110111011101111111111101111111111101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101110111011101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111101110111011111111111111111111111011101110111011101110111011101110111011011101110011001100101111001100110011001100101111001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011100100110010001000100101101010111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110001001100010001000100010001000100010000100001000100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100001001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000110100010001000011001100110011001100110010001000100011001100100010001000100010001000100010001100100010001100110011001000100010001000110011001100110011010001000100001100110100011110111100110011001101110111011101110111011101110111011101110111011101110111011101110111011100110011011100110110110111010000110100010000110011001101000100010001000100001100110100011110011000010101000100010101110111010101010101010101000011001101000011001100110100010000110010001000110101010000110011001100110011001101000100010001000101011001110111011101100110011001010101010101101000100110111100110111011100100110000101010001111110111011101110111011101110111011101110111011101110011101111110111011101110111010010111111011101110111011111111111011101111111111111111111111111111101010001110111111101110100010111110110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101111111011111111111111111111111011101110110111011100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011100101000010001000100101101010111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010000101001000100010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110010001000100010001000100010001000100010001000100010001100100011001100110011001100110011001100110011001100110011001100110100100010111100110011001101110111011101110111011101110111011101110111011101110111011101110111011100110111011101110110010100010001000100010000110011010001000100010001000011001101000111101010101000010001000101011001100110010101100110010101000100010001000011001100110100010001000010001000110101010000110011001100110011010001000100010001000100010101100111011101100110011001100101011001010110011110001001101111011100100110000101010010011110111011101111111011111110111111101110111011111110011010011110111011101110111010001000111011101110111011111111111011101111111111111111111111111110100010101110111011111100011111011110110111011110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011111111111111101110110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011100101000010001000100100101010111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010000110001000010010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001000100011001101000011001100110011001100100010001000100010001000100010001000100010001000100010001000100011001100100011001100110011001100110011001101000100011110111100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101101110101010001000101010100110100010001010101010101000011001101011001101110100111010001000110011101100111011101110110010101010100010001000011001100110100010001000010001001000100010000110011001100110011010001000100010101000100010101100110011001100111011001100111011101100110011001110111011110011001100101110100010010111110111011101111111111111111111111111111111011111100010110111111111011101111110101111010111111111111111011101111111111111111111111111111111111111100011110111111111111111001100011101110111011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111110110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101001000010001000100100100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010000110001000010010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000010001001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110100010001000100010110001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100101100101010001000110011001000100011001111000010101000100010010001011110010100110010001010111011101111000100010000111011001010101010101000011001100110101010101000011001001000101010000110011001100110011010001010101010101010101010101010110011110001000100001111000100001111000011101100110011001100111100101100100011011011110111011101111111111111110111111111110111011111011010111011111111111101111110001101100111111111111111111111111111111111111111111111111111111111010011111011110111011011000101111111110111111101110111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001000010001000100011100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010000111001100100010001000110011010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100100010001000100001001000100010001000100010001000100010001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001010101010101010111110011011101110111011101110111011101110111011101110111011101110111011110111011101110110111011011100001100101010101010111011001000100100010101000010101000100010110111100101110010101010101111000100010001001100010001000011001100110011001000100001101000101010101000011001001000100010000110011001100110011010001010101010101010110010101010110011110001001101010001001101010011000100101110110011001100110011101010100100011101111111011101111111111111110111111111110111011111001011111101111111111101111101101101101111111111111111111111111111011101110110111011101110011001000100011011101111010111000110111101110111011101110111111101111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001010010001000100011100010111011101110111011101110111011101110111011101110111010101110111011101110111011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000001100010010001000110011010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001010101010101010100011110111101110111011101110111011101110111011101110111011101111011101110111011101110110111001010100101110110011001101001011101000101101010111001011001000100100011001100101101100100011010001001100110011001100110011001011101110111011001000100010001010101010101000011001101000100010000110011001100110011010001010101010101010110011001010101011001111001101010101010101010111001101010011001011101100110100001010101101011101110111111111111111111111111111111111111111111100111100011101111111111101111101001111110111111101111111111111101110010111011101110101010101010010111100110101011101110011001110011011110111011011110111111101110111011101111111011111111111111111111111111101101110111011110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001010010001000100010011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000010000010001001000010010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000010001000100100010001000100010001000100010001000100010001000100011001100110100010001000100010101000100010001101010110111011101110111011101110111011101110111011101110111101110111011101110110111001011101010011000011110001010011101000110101111001010010101000110101111011100100101010100011110011001100110011001100110101010100110011000011001000100010001010101010101000011001101010100010001000100001100110011001101000110011001100111011101100110011001111000100110101010101111001011101010111011100101100111011101000110110011111110111111111111111111111111111111111111111111010110101011101110111011101110100010001110111111111111111011011100101110101010101010101010101010010111100110011001100110001001101010111100110011011110111011101110111011101110111011101111111111111110110111011101110111011101110111011101111011011101111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001010010001000100010011010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000010100010001001000100010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100010001001000100010001000100010001000100010001000100011001100110011001101000100010001000100010001000111110011011101110111011101110111011101110111011101111011101110111011101101110111011100110011001010100110011100011101010111110011000111010001001001110111001011011101010101100110101010101010101010101010111011101110101000011101010100010001010110011101100011001101010100010001000100001100110011010001000110011001100111100001110111011101110111100010011001101010111100101010111100101110101001011001000111111011111111111111111111111111111111111111111111111111000110110011101110111011101100011010101111111111111101101110101010101010101010101010101010101010000111100110011001100010001001100110011010101010111100110011011110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101001100010001000100010010110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100010001000100010001000100010001000011000100001000100010010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001000100100011001100110010001000100010001000100010001100110011001100110100010001000100011010011100110111011101110111011101110111011101110111101110111011101110111011101101110111011101111011011100101110111101011101011000110010100101010001101100110111001001011001010111100110101010101010101011101111001100101110101001011101010100010101111001101001110011010001010100010001010100001100110011010001000101011101110111011110001000100010001001101010101011101110111100101110011011110011001010010101001010111011111111111111111111111111111111111111111111111110100110110111101110111011101010011010111101110010111010101010101010101010101010101010101010100101111000100110011001100010001001100110011001100110011010101010101011101111001100110111011101110010111100110011001101110111011101110111011101110111011101110111011101110111011110111011111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001110010001000100010010110101011101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000011100100001000100100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001100110011001100110100010001011000101111011101110111011101110111011101110111011101110111101110111011101110111011101101111011101110111011101101110011011101011101011000101101110101010110101101110110110111010101011000101010101010101010101011101111001100101010011000011001000100011110111101110001110011010001100110011001100100001100110011010001000110100110011000100010001001100110111100110011011101110111011101110010101010110011001001010001101100111111111111111111111111111111111111111111111111111110010111110011001100101110110111011010101010101010011001101010101010101010101010101010101010100101111000100110011001100010011001100110011001100110011001100110011001100110101010101010101010100110011010101010101010101110111100110011011101110111011101110111011101110111011101111011101110111011101110110111011101110111011110111011101111111111111111111111111110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001110010001000100010010010101011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100010001001100000110001000100010010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010010001000100010000100100010001000100010001000110011001101000101010101101000110011011101110111011101110111011101110111011101110111011101110111101101110111011101111011101110111011101110111011101101011001010110011101010101011111011101110010010101010001101010101010101010101010101010101010111010101010010111010101000101100010111100101101100011011010011000011101010100001100110011010001000111101110101011101010101100101111011101111011101110111011101110110111001010110011000111010001111110111111111111111111111111111111111111111111111111111001110110100110011000100110000101011110011001100110011001101010101010101010101010101010011001100001111001100110011000100010011001100110011001100110011001100110011001100110011001101010011001100110011001100110011001100110101010101010101011110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011111111111111111111111111111111111011101111111111111111111111111111111111111111111111011100110111011110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010000010001000100010001110011011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100000110001000100010001001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100011001101000100010001011000110011011101110111011101110111011101110111011101110010111011110111101110110111101110111011101110111011101110111011101100011001010101010101010110101111011101101101100101010010001011110010111011101010101001100110011010101010000111010101000100011110111101110110000011100010101001011001000100001100110100010001000111110011001100110011011101110111101110111011101110111011101110111011011010101010110101010010011110111111111111111111111111111111111111111111111111110101010111100010001000100101110101011110011001100110011001100110011001101010011010101010011001100001111001100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110011010101010111011110011001101110111011101110111011101110111001100110111011101110011001101110111011101110111011101110111011101110111011101110111101110111011101110111011101110110111011110111011101110111011101110111011101110110111011101110111011110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010000010001000100010001110001011101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100001000001000100010010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001100110011010110001100110111011101110111011100110011001011101110101001100001111000110011011101110111011110111011101110111011101110111011101100011001010101010101011000110111001100100001010100010110101101111011001011101010011001101010101011101010010111010101000100100111001101110101110011100010100111010101000100001100110011010001000111110011011101110111101110111011101110111011101110111011101110111011001011101010010100010110111111111111111111111111111111111111111111111111111111101001011000100010001001100001100101100010011001100110011001100110011001100110011001100110011001011110001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011010101010111100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110010011001000100001001010001011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100001010001000100010010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001100110100011110111101110110111010100110010111011101110110010101010100010000110101100011001101110111011110111011101110111011101110111011101010010101010101010101111100110010111001010101000100011110111101111011011011101010101010101010111011100110000111010101000101100010111100101101100011100010010111010101000100010000110011010001000111110011001100110111101110111011101110111011101110111011101101101110101011101001110100011111011111111111111111111111111111111111111111111111111110011101011001100110011001100001010110100010011001100110011001100110011001100110011001100110011001011110001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010111011101110111011101110111011101110111011101111001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010010011001000100010001001111011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100101100010000100010010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000110011001101000101011110001000011001010100001101000100010001000100001100110011001100110101100111001101111011101110111011101110111011101110111011101001010101010110011110101100101010010111010001000101100110111011101110111010100110011010101110111001100110000110010101000101100010011011101101010100100110010110010001000100001100110011010001000110101010111011110011011110111011101110111011011100110011001100101010001001100101010100100011101111111111111111111111111111111111111111111111101100010101101001100110011001011101000110100110011001100110011001100110011001100110011001100110011000011110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101011101110111011110011001100110010111011101111001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010100100001000100010001001111011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100101110010001000100010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001100110011001101000100010000110011001100110011001100110011001100110011001100110011001101000101011110011100110111011110111011101110111011101110111011101000010101010110101010111011100110000101010001000110100010001000100010001000100001111000100010001000011101110110010101000101011110001001100101000011011110000110010001000100001100110011010001000101100010001000100110111100110011001100110010111010100110001000100010001001011101000100101011111111111111111111111111111111111111111111111011011010010010001001100110011000011001000111100110011001100110011001100110011001100110011001100110010111011110011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101111001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010100100001000100010001001101011101110101011101110111011101010111010101010111011101010101011101110111010101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010000100001000010010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001000100001000100010001000100100010000100010001000100010010001000100010001000100010001100110011001100110010001000100010001100110011001100110011001100110011010000110011001100110011001101000110100010101100110111101110111011101110111011010111010101010111110010101001100101100100001101000110011101110111011101110111011101100111011101110111011101100101010101000101011101111000011101000011011001100101010000110011001100110100010001000100011001110110011101111000100010001001100110011001100001110111011110001001011000110101101111101110111111111111111111111111111111111110110111011001010110011001100110011000010101011000100110011001100110011001100110011001100110011001100110010111100010011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101111001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010100101001000100010001001011010101110101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000100000100010001001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001001000010001001000100010001000100010001000100010001000100010001100110011001100110011001100110100001100110011001100110011001100110011001101000110100010101100110111101110110110110110010001011001101110011001011101000011001101010111011101110111011101110111011001100110011001110111011001100101010001000101011001110111011000110011010101010100010001000100001100110100010101010100011001100110011001100110011001110111011101111000100010000111011101110111010000110110101011001101110011011110111111111110110111001101111011101000010110011001100010000111010001101001100110011001100110011001100110011001100110011001100110000110100010011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101111001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010100110001000100010001001011010101110101011101110101010101010101011101010111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000101001000010010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100100010001000100001000100010001001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110100001100110011001100110011001100110011001100110011001101000110100111001100110010100101010001011001101010101000010101000011010001100111011001100110011101110111011001100110011001110111011001100101010001010101011001100110011000110011010101010101010001000100010001000100010101010101011001100110011001100110011001100110011001110111100001110110011001100110010000110110011110011010100010011100111011111101101110111101111011010110011010000111011001110110001101111001100110011001100110011001100110011001100110011001100101110110100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101111001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010100111001000100010001001001010101110111011101010101010101010101010101110111010101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000110001000010001001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001100110011001100110010001000100011001100110011001100110011001100110100011010011010101110010100010001001001101010010111010000110011010001100111011001100111011101110111011001100110011101100111011001100101010001010110011001100111011000110100010101100110010101000100010001000100010101100101011001100110011001100110011001100110011001100111011101110110010101010100001101000101011001111000011101111001110111011010011110001000101010010100011001110101010101010100010010001001100110011001100110011001100110001000100110011001100101110111100110011001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010100111001000100010001101001001101110101010101010101010101010101010101010111010101010111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010010111001000010010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000010001001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001000100010001000100011001100110011010001000100010101111000100101110100001101001000100110010101001100110011010001100111011101110111011101110111011001100111011001110110011101100101010101010110011001110110010100110100011001100110010101000100010001000100010101100101010101100110011001100110011001100110011001100110011001100101010101010100001101000101010101100111011001110111101110010110011001100110011001010100010101100101010101010100010110001001100110011001100110011001100101110111100110011001100001101000100110011001100001111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101111001100110011001100110011001101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010100111001000100010001101001001101110101010101010101010101010101010101010101010101110101010101010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000001100010010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010000100010001001000010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001000100010001000100010001100110011010001000100010101110111011101010011001101011001100101110011010001000100010001100111011101110111011101110111011001100110011001100110011001100101010101100110011001100110010100110101011001100110011001010101010001000101011001100110010101100110011001100110011001100110010101010101010101010101010001000011001101000101010101010110011001100110011101100101010101010101010101010100010001010101011001010011010101110111100010011000100010001001100101110110011110001001011101101000100010000111011001111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011110011001100110011001100110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101000001100100010001000111000101110101010101010101010101010101010101010101010101010101010101010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010000100010001000100001001001101000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100001001000010001000100100001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001010110011001000011001101101001100101010011010000110011010101100111011101110111011101100110011001100110011001100110011001010100010101100110011001100110010000110101011001100110011001010101010101000101011001100110010101100110011001100110011001010101010101010101010101010100010001000011001101000101010101010101011001100110011001100101010101010101010101000100010001000100010101000011010101100110011101110111011110001001100101110101011001111000011001100111011101100110010101100111100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011110011001100110011001100110011001101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101000001100100010001000101000101110101010101010101010101010101010101010101010101010101010101010111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010100100010001000100001000101011000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000010001001000010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010000110010001101011000011000110100010000110011010101100110011001100110011001100110011001100110011001100110011001010100010101100110011001100110010000110110011001100110011001100110010101010101011001100110010101010101010101010101010101010101010101010101010001000100010001000011010001000101010101010101011001100110011001010101010101010101010101000100010001000100010000110100010101010101011001100110011001100111100001110110011001100110010101100111011101100101010101010110011101111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111100110011001100110011001100110011011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101001001100100010001000100111101110101010101010101010101010101010101010101010101010101010101010111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001101010101001100110101001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011000100010001000100001000101001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000110010001100110011001100110011001101010111010001000100001100110100010101100110011001100110011001100110011001100110011001100110011001010101010101100110011001100101010000110110011001100110011001100110011001010110011001100101010101010101010101000100010001000101010101010100010001000100010000110011010001000101010101010101011001100110011001010101010101010101010001000100010001000100010000110100010101010101010101100110011001100110011101110110011001110101010101111000011101010100010001000101010101100111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011110011001100110011001100110011001100110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101001001100100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100100010001000100001000100110111100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100100011001101100110010001000011001100110100010101010101011001100110011001100110011001100110011001100110010101000101010101010100010101010101001101000110011001100110011001100110011001100110010101010101010101010101010101000100010001000101010101010100010001000100010000110011010001000100010001000101010101100110010101010101010101010101010001000100010001000100010000110100010101010101010101010110011001100110011001100110010101010100010101100101010101000100010001000100010101010111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101011101010111011101111001100110011001100110011001100110011001100110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011110010111100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101001010000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100110010001000100001000100100111100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100010001001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100100010001101010101010001000011001100110100010101010110011001100110011001100110011001100110011001100110010001000100010001000100010001000100001101000110011001100110011001100110011001100101010101010100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000101010101010101010101010101010101010100010001000100010001000100001100110100010101010101011001010101010101010110010101010100010001000100010001000100010001000100010001000100010001010110011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111100110011001100110011001100110011001100110011001101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101001010000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100000110001001000100001000100100110100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000010010001000010001000100010001000100010001000100010001001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000010001001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010101010100001100100010001101010101011000110011001100110100010101010101010101100110011001100110011001100110011001010100001100110100010001000100010001000011001101000101010101100110011001100110011001010101010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000100010001000101010101010100010101010100010001000100010001000100001101000100010101010101011001100101010101100110010101010100010000110100010001000011010001000100010001000100010001010110011110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101100111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001100010011010101010101010101010101010101010101010101010101010101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010010000100010001000100101101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100001000010001000100001000100010101100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000010010000100010010000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000110100010101010101001000100011010001100111011000110011001100110100010101010101010101010101010101000100010001010110011001010100001101000101010101010101010101010011001101000101010101010101010101100110010101010100010001000100010001000100010001000100010001000100010101010100010001000100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001101000100010001010101010101100101010101010110010101010100001101000100010001000011001100110100010001000100010101010110011101111000100010001001100110011001100110011001100110011001100110011001100010001001100110011001100001111001100110010111011001010110011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001100010011010101010101010101010101010101010101010101010101010101010111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100101110111100110011001100110010111011101110111011101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010010100100010001000100101101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010001000100010000100010100100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000010010001000010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000110011001100110100010101010011001000110011011001100101010000110011001100110100010101010101010101000100010001000100010001010110011001010011001101000101010101010100010001000011001101000101010101010101010101010101010101010100010001000100010001000100010001000100010001010100010001000100010001000100001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001101000100010001000101010101010101010101010101010101000100001100110100010001000011001100110011010001000100010101100110011101110111011110001000100010001001100110001000100110011001100110011001100001111000100110011001100001111000100110000111011001100111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111100010011001100010001000100010001001101010101010101010101010101010101010101010101010101010111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010011000100010001000100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100010001000010011011110001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001100110100010101000010001000110011011101100100001100110011001100110100010001000100010001000100010001000101011001100110010101000011010001010100010001000100010001000011001101000101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010000110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010101010101010101010101010001000011010000110100010001000011001100110011010001000100010101010101011001100111011110001000100010001000100010001000100010001000100010011000100001111000100110011001100001111000100110000110011001100111100010011001100110011001100110011001100110011001100110011001100110011001100110000111100001100110011110001000100001110111011001100111100110101010101010101010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111010011000100010001000100100101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110010001000100010001000010010011010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100100011001000100010001000100010001000100010001000100010001000100010000100100001001000100010000100100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100100010001000100011001100110010001100100011010101110100001100110011001101000100001100110100010001000100010001010110011001100110010100110011010001000100010001000100010001000011001101000101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010000110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010101010101010101010101010001000100010000110011010001000100001100110011010001000100010101010101010001010110011110001000100010001000100010001000100010001000100010001000100001110111100010001000100001111000100001110111011001100111100010011001100110011001100110011001100110011001100110011001100110011001100101110111011001010101011110000111011101110110010101010110100110011010101010101010101010101010101010101010101010101010101110111011101110101010101010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010011100100010001000100011100110111010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000011000100100001000100010010010110001000100010001000100010001000100010001000100010001000100010001000,
	2400'b010101010101010101100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001000100010001000100010001100100011010101110100001100110011001100110011001100110100010001000100010101010110011001100110010000110011010001000100010001000100010001000011001101000100010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010101010101010101010100010001000011010001000011010001000100001100110011010001000100010001000101010001010101011001111000100010001000100010001000100010001000100010001000100001110110011101111000100010000111011101110111011001100110011110001000100010001000100110011001100010001000100010001001100110011001100001110110011001010101011010000111011101100101010101010110011110001001100110011001100110011001101010101010101010101010101010111011101010001000100010101011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100100010001000010011100110111010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100010001010010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b010101100101010101100101001101000101010000110010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110010001000100010001100100011010001010011001100110011001100110011010001000011001100110100010101010110011001100101010000110100010001000100010001000100010000110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010001000100010001000100010001000100010001000011001100110100010001000100010001000100010101010101011001110111011110001000100010001000100010001000100001110111011101110110011001100111011101110111011101110110011101100110011110001000011101100111100010011000011101110111011001101000100110011001100001110110011001010101011001100111011101100101010101100110011001111000100010001000100010011001100110011001101010101010101010111010101010001000100010011010101010101011101110111011110011001100101111001100110011001100101110101001101111001100110010111100101111001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100000100010001000010010100010111010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101110111011101010101010101010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010001000100010001001110001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100110011010001000011001101000101010101010100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001000100011001000100011010001000011001100110011001100110011001101000011001100110100010001000101010101010100001100110100010001000100010001000100010000110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010000110011001100110100010001000100010101000100010001010101011001110111011001100110011110001000100001111000100001110110011001100110011001010110011001100110011001100110011101100110011101110111011101100110011110001000011101100110011001101000100110011001100001100110011001010101010101100110100001110110011001100110011001110111011101110111100010001001100110011000100110011010101010101010101010010111011101111000100010001010101110111011101110101001100110101011101111001011100101110110100010111100110011001100101110111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100100110010001000100010011110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000010001000100010001001001111001100110001001100110011000100110011001100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001000100011001000100011001100110011001100110011001101000011001100110011001100110011010001000100010001000100001100110100010001000011010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010001000100010001000100010001000100010000110100010001000100010001000011001100110011010001000101010101010101010101010101011001110110010101010101011010001000011101110111011001100110011001010101011001010101011001100110011001100110011101100110011101110111011101100110011001111000011101100110011001101000100010001000100001100110011001010101011001100110100010000111011001100110011001110111011101110111011101111000100010011000100010001001100110101010101010011000011101110111011101111001101110111011101001110110011110011010101111001011100001100110011110101100110011001100101010001000100010111011101110111011101110111011101110111011101110111011101110111011110010111011101111001011101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000110010001000100010011110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000010001000100010001001001101001100110011001100110011001100010011001100010011000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110010001000110010001000100011001100110011001100110011001101000100001100110011001100110100010001000100010001000011001101000100010001000100010001000100001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011010001000101010101010101010101010101011001100101010001010101011001110111011101110110011001100110011001010101010101010101011001100110011001100110011101110111011101110111011101100110011001111000011101100110011001110111011110001000100010001000011101100110011001100111100010000111011001100110011001110110011101110111011101110111011110001000011101110111011110001001100110011000011101100110011001111001101110111001100001100110011110011001101110111011100001100111100110111100110011001011100101110111100010111011101110101010101010111011101110111011101110111011101110111100110010111011110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101001000010001000100010011010111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111001000010001000100010001001001011001100110011001100110011001100110011000100110011001100010011000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110010001000110010001000110011001100110011001100110011001100110100010000110011001100110100010001000100010000110011001101000100010001000100010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000101010101010101010101000100010101100101010101010101011001100101010101100110011001010101010101010101010101010101011001100110011001100110011001100110011101110111011101100110011001100111011101100110011101110110011001110111100010000111011001100110011001100111100010000111011001100110011001110110011001110111011101110111011101111000011101100110011101110111011110001000011101100111011001111010101110101000011101100110011001111000101110111010100101111001110011001100110010111011100110000111011110111011101110000111100010101011101110111011101110111011101110111011101111001011101111001100110011001100110011001100110010111011101110111011101110111011101110111011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101001010010001000100010010110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000001100010001000100010001000101001000100110011001100110011001100110011001100110011001100110011000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100100010001000100010001000110011001100110011001100110011001100110011001100110011001100110100010001000100010000110011001101000100010001000100010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010101010101010001000100010001010101010001010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110011001100111100010000111011001100101011001100110011001100110011001110111011101110111011001100110011001100110011001100111011001111000100010011001100110101000011101110110011001110111100110011001100001111000101110111100110010111010101010010111011110011011100101110111011110011011101110111011101110101010101110011000101111001100110011001100110010111011110011001100110011001100110010111100110011001011101110111100101110111011101110111100101110111100110011001011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101101010010001000100010010110101011101010101010101110101010101010101010101010101010101010101011101110101011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010000100001000100010001000100111000100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100100010001000100010001000110011001100110011001100110011001100110011001100110011001100110100010001000100010000110011010001000100010001000100010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001101000100010001000100010001000100010001000100010001000100010101010100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101011001100110011001010110011001100110010101100101011001100110010101010110011001100110011001100110011001100110011001110111011101110111011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011110001000011101110110011001110110100010010111011101110111100010101011101110111001101010000111011110001010101010000111011110001011101110111011101110001000100101100111101110101001100110101011101111001100110011001100110011001100101110101011101110111011110010111100101110111100110011001100110011001100101110111011110011001100101110111011101110111011101110111011101110111011101110111011101110111011101101100010001000100001010010101011101010101011101110101010101010101010101010101010101010111010101010111011101110111011101110111011101110111011101110111011101110111010101110111010101010111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010100110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010000010001000100010010000100100111100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001100110011001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110100010001000100001100110011010001000100010001000100010000110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100111011101110110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101111000101011001010011101110111011110001010101010011000100010001010101110111011101010001000011101010110100001110110011001111000101011001100110010111001100110101011101010011001100110101011101110111011110011001100110011001100110011001100110010111100110011001011101110111100110011001011101110111011101110111011101110111011101110111011101101110010001000100010001110101011101110111011101110111010101010101010101110111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010101010101010101010100110101010101010101010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100100001000100010001000100100110100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001100110011001000100010001000100010001100110011001100110011001100110011001100110011001100110011001101000100010001000100001100110100010001000100010001000100010000110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111100001110111011101110111011101110111011101110111100010011000011101110111011110001001100010001000100010011010101010111011101010010111011001100110011001100111011001110111100110111010101010010111011110001001100110001000100010011001100110101010101110111010101010101010101110111011101111001011101110111011101111001100110011001100110010111100110010111011101110111011101110111011101110000010001000100001001110011011101110111011101110111010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011000100001000100010001000100100101100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000110011001000100011001000100010001100110011001100110010001100110011001100110011001100110011001100110100010001000100001100110100010001000100010001000100010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101111000011110000111100010001000100010011000100010001000100110101001011101100110011001110111011101111001100110011000100010000111011101110111100010001000100010001000100010001000100010000111011101110111011110001001101010101010101010111011101110111011101110111100110011001100110011001011101110111011101110111011101110000010001000100010001010011011101110111011101010101010101110101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101010101010101010101010101010101010101010101010011010100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100100001000100010001000100010100100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100100010001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000110011001100110011001000100010001000100010001000100011001000100010001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010000110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110100010001000100010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001001011110000111011101110111011110000111011101110111100110111001100001110111100001110111011101111000100010001000011101111000100010001000100010001000100010001000100010000111011101110111011101110111011110001000100010001000100110011010101110111011101010011011110011001100110011001100110010111011101110111011110010010010001000100010001010001011101110111010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100000110010000100010001000100010011100010011001100110011001100110011001100110011001100110011001,
	2400'b001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100100010001000100010001100110011001000100011001100110011001100110011001100100010001000100010001000110011001100110011001000100010001000100010001000100011001000100010001100110011001100110011001100110011001100110011001100110011001100110010001000100010001100110011001101000100010001000100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000101010101010101010101010101010101010101010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010000111011101110111011101110111011101111000101010101000100010001000100101110111011101111000100010001000011101111000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001001100110101011101110111011110011001100110011001100110011001011110010111011110010010011001000100010001001111011101110101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010111010101110111011101110111010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010001000010010001000010011100010011001100110011001100110011001100110011001100110011001,
	2400'b010001000100010000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100100010001000100010001100110011001000110011010001000100010000110011001100110011001000100010001000110011001100110011001000100010001000100010001000110011001000100011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001000100010001100110011001101000100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010001010101010101010101010101010101010101010101010101010101010101000101010101010101010101010101010101010101010101101000100001110110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101111000100010000111011110001000100010001000100010001000100010001000100001111000100010001000100001111000100110001000100010001000100110000111011110001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011010101111001100110011001100110011001100110011001100110011001100110010010011000100100010001001101011101110101010101010111010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010001000100010001000100010011110011001100110011001100110011001100110011001100110011001,
	2400'b010000110011001101000100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100100010001000100011001100110011001100110011010001000100010000110011001100110011001000100010001000110011001100110011001100100010001000100010001000110010001000100011001100110011001100110011001100110100010001000100010001000100010000110011001100110011001100110011001100110011001100110100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010101010101100110010101010101010101010111011101100110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001101010111011101110111100110011001100110011001100110011001100110010010010001000100010001001001010101110111010101010101011101010101011101010111010101110111011101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101110111010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010011001101010011001100110011001100110011001100110011001100110011001100110011001100101100010001000100010001000100010011010011001100110011001100110011001100110011001100110011001,
	2400'b001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001000100011001100110011001100110100010101010101010000110011001100110011001000100010001100110011001100110011001100100010001000100010001100110010001000110011001100110011001100100011001100110100010001000101010001000100010001000100010001000011001100110011001101000011001101000011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010101011001100111011001010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011010101010101011101110111011110011001100110011001100110010010011000100100010001000111010101110111010101010101010101010111011101010101011101110111011101110101010101010101011101110111011101110111011101110111100101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110101010101010101010100110011001100110011001100110011010100110101010101010101010101010101010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101001110010001000100010001000100010010110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100100011001100110011001101000100010101010101010000110011001100110011001000100010001100110011001100110011001100100010001000100010001100110010001100110011001100110011001100110011001100110100010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000100010001010110011001100101010001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011101010101010101100110011010001000011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011010101010101010101111001100110011001100110010100011001000100010001000111010101110111010101010111010101010101010101010111011101110111011101010011010101010101011101110111011101110111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101010011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001101010000011001000100010001000100001010010011001100110011001100110011001100110011001100110011001,
	2400'b001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100100011001000100010001000100011001100110011001000100010001000100011001100100010001000100010001000110011001100110011001100110011001100110011001100110011001101000101010101100110010001000100001100110011001000100010001100110011001100110011001000100010001000100010001100110010001100110011001100110011001100110011001100110101011110001000100110001000011101100101010101010100010001000100010001000100010000110100011001110111011101110110010101000011001100110100010001000100010001000100010001000100010001000100010001000100001100110011001100110100010001000100010001000100010001000100010001010100010001000011010001011000101010000101011001100101010101000100010101000100010001000100010001000100001101000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100101011001100110011001111000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011110001000011101110111011110001000100010001000100010001000100010001000100010001001100010001000100010011001100110011001100110011000100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101110111011101110101010101010010011001000100010001000111001101110111010101110111010101010111010101010111011101110111011101010101010101110111011101110111011101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010100110011001100110011001100110011001101010101001100110011001100110011010100110011001100110101010100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010100110101010100110011001100110011001100110101010101010101001101010010011001000100001000100010001001110001001100110011001100110011001100110011001100110011001,
	2400'b001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100100011001100110011001000110011001100110011001100100010001000110011001100100010001000100010001100110011001100110011001100110011001100110011001101000011001101000101010101010101010010000111001100110011001000100011001100110011001100110011001000100010001000100010001100110011001100110011001100110010001100110011001101000110011110001001100110011001100110000111010101010100010001000100010001000100010101010100010110011100100101110111100001100011001100110100010101000100010001000100010001000100010001000100010001000011001100110011001100110100010001000100010001000100010001000100010001000100010000110011001101010110100001110101011001100111011001010100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001010101011001100111011001100101010101010101010101010101011001100110011001100110011001100110010101100101010101100110011110001010101010101000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100101110111011101110111011101110111011101110111011101110111011101110111011110001000100010000111011101111000100010001000100010001000100010001000100010001000100010011000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101001100110011001100110010011000100100010001000101000101110101010101010101010101010101010101010101010101010101010101010101010101010111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100000100100010000100010001001110001001100110011001100110011001100110011001100110011001,
	2400'b010001000011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000110010001100110011001100110011001100110011001100110010001100110011001100110010001000100011001100110011001100110011001100110011001100110011001100110100010001000100010001000100001110001000001100110010001000100011001100110011001100110011001000100010001000100010001000100011001100110011001100100010001100110011001100110101011101111000100110011001100001110111010101000100010001000100010001000100100110010100010010011100100001010101100001110100010000110100010101000100010001000100010001000100010001000100010001000100010001000100010101010100011001100100010001100111011101100110010101010101010101010100010110000110010101010101010101100111100110000110010101000100010001000011001100110011001101000100010001000100010001000100010001000100010001010101010101100111100010001000100010000110011001100110011001100110011001110111011101110111100010000110010101100111100010000111011101111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010000111100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011010100110101001101010101010101010101010101010101010101010101010100110101001101010101010100110011001100110011010100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001100110011001100110010100000100100010001000100111101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110110110001000100010001000010010001010001010101010101010101010101010101010101010101010101010,
	2400'b100001110110001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001100110011001100110011001100110011001100110011001100110011001100100011001000100011001100110011001100110011001100110011001100110100010000110100010100110011001100110011001100110011001100110011001000110011001100110011001100110011001000100010001000100010001000100010001100110011001100100010001000110011001100110100011010001000100010001000100001110110010001000100010001000100010001000100100110100101010010001010100001000101011101110100010000110011001100110011001101000100010001000101010101010110010101010101011001100110100010010111101010100110001101111001100110011001100110001001101010011000100110101000011001010101010001000100010101010110010101000011001100110011001100110011001101000100010001010101010101000100010001000101011001110111100010011001100110011001100110101001100010001001100110011001100110011010101010101011101110111010011110011101111011011010101010101010101110111010101010101001100110001000100010001000100010001000100010001000100010001000100110101001100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110001000100110011001100110011001100110011001101010101010101010101010101010101011101110111011101110111011101110111011101111001100101111001100110011001100101110111011101110101010101010111011101110111010101010101010101010101011101010111011101110111011101010101010101110111011101110111011101010101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010010100000100100010001000100110101010101010101010111010101010111011101110111011101110111011101110111011101110111100101110111011101110111100101110111011101110111011101110111011110010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011110011001000001000100010001000100010001001111100110011001100110011001100110011001100110011001100,
	2400'b100110000111001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100100010001000110011001100110011001100110011001101000100010001000100010000110100001100100010001100100010001100110011001100110011001000110011001100110011001100110010001000100010001000100010001000100010001100110011001100110010001000110011001100110011010101111000100010001000011101100101010001000011001100110011010000110100010101100100010001101000011001000101011001100100001100110011001100110011001100110100010001000101011001110111011101100110011101111000100010000111100110010111010101010111011001100111011101110111011101110110011001100101010101010101010001000100010001000100010001000011001101000011001100110011001101000100010101010101010001000100010101111001101010111011101110111100101110111011110011001100110010101011110011001100110011001100110111011101110111011100011110001100110011001100110011001100110011001100110011001100101110101010101010101010101110111011101110111011101110111010101111001101101110101100110011001100110011001100110011001100110011001100110111011101110111011101110111001100110011001100110011001100110011001100110011001100110111011101110111011100110011011100110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110111001011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111100101110111011101110111100110011001100110011001100110011001100110011001100110010111011101110111011101110110101000100100010001000100110101110111011110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101101110111011101110111101110110111011101110111011101111011101110111011101110111011101110110111101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001101110111011100110011011101110011001100110011001100110011001100110011001100110011001100110011011001001000100010001000010010001001101101110111011101110111011101110111001100110011001100,
	2400'b100110000111001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100100010001100100010001100100011001100110011001100110011001100110011001000100010001000110011001100110011001100110011010101010110011001010100010000110011001100110011001100110011001100100011001100110011001100110011001100110011001100110010001000100010001000100010001000100010001100110011001100100010001000110011001100110011010001100110011001100110011001010100010000110011001100110011001101000011001101000100010001000100010001000100010001000100001100110011001101000011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101000101010001000100010001000100010001000100010001010101010101100101010101100110011010001010110011001100110011001100110011001100110111011100110111011101110011011101110111011101110111011101110111011101100010011011110011001101110111011100110011001101110111001100110011001011101111001100110111011101110111011101110111001011101111001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011100110011001011110011001100110011001100110011001100110011001100110011001100110011001100110111011101110011001101110111011101110111011101110111011101110111001011110011001100110011001100110011001011101110111011101110111011101110111011101110111100110011001100110011001101110011001100110011000111000100100010001000100110110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011010001100100010001000010010001001011100110111011101110111011101110111011101110111011101,
	2400'b011001010100001100100010001000100010001000100010001000100010001000110011001100110011001000100010001000100010001100110010001000100010001000100010001000110011001100110011001100110011001000100010001000100010001100110011001100110011001100110100011110000111011001010100001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001000100010001000100010001000100011001100110011001100110010001100110011001100110011001100110100010001000100010101000100010001000100010001000100010001000100010001000100010001010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010110011101111000100010011001100110011001100110101010101111001100110011001100110111001100110011001100110111001101110011001100110011011101110111011101110111011100101010101100110011001100110011001100110011001100110111011101110111011100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111001100110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110011001100110011001101110111001100110011001011101110111100110011001100110011011101110011001100110011001100110011011100110011011101111011101110111011101110111011101110111011111001000100100010001000010101111011101110111011101110111011101110111011101110111111101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111101110110111101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011010000100010001000010001001000111011110111011101110111011101110111011101110111011101,
	2400'b001100110011001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001100100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011010001000100010101010110011001010101010001000011001100110011001100110100010001000100010001010100010101010100001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001101000100010001000100010001000101010101010101010101010101010101010100010001000100010101010101010101010110011001100111011101100110010101000100010101010101011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101000100110011010101010101010101010101011101110111011110011001100110011001100110011001101110111001101110111011100110011001101110011001100110011001100110011011101110010111100100110011100110011011101110111011101110111011101110111011101110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001101110011001101110111011101110111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011011110111011101110111011011110111011101110111011101110111011101110111011101110111011101110110111101111111111101110111011101110111011101110111011111010001000100010001000010101111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111101110110111011101111011101110110111101110111011011101110111011101110111011101110111011101110111011101110111011100010100100010000100010001001000111001110111011101110111011101110111011101110111011101,
	2400'b001100110011001100110011001100110011001100110011001100110011001101000100010001000011001100110011001100110011001100110010001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010101010101010101010100010001000100010000110011001100110011010001000100010101010101011001100100010001000100010101000110011001000011001100110011001100110011001100110011001100110011001100110011001101000100010001010101010101010101010101010101010101010101010101000100010001000100010001010101010101010101010101010101011001010101010101000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011101110110011001100110011001100110011001100111100010001001100110011001101010101010101110111100110011001100110111011100110011001101110111011100110011001100110010111011101110111011101110111011101110111011101110111011100110101100110111011101110111011101110111011101110111011101110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100101111001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110110111101110111011101110111011101110111011101110111011101110111011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011111100001100010010001000100100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101101110111011101110111011101110111011101011000100001000100100010001000101000110111011101110111011101110111011101110111011101,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011001100110011001100110011010001000100010101010101010101000100010001000100010000110011001100110011001100110011001100110011001101000100010001000100010001010100010001010101010101010101010101000100010001000100010001010101010101010101010101010101010101010101010001000100010001000100010001000100010101000100010001000101010001000100010001000101010101010100010101010101010101010101010101010101010101010110011001100110011101110111011110000111100001110111011101110111011101110111011101110111011001100110011001100110011001110111011101111000100010001001100110101010101010111011110011001100110011001100110011001100101110111010101010011001100110011001100110011001100110011001101010101010101111001100110011001100110011001100110011001100110011001100110011001100110111011100110011001101110111011101110011001100110011001100110011011100110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111101110111011101110111011111110111111111110111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111011111111111011111101001100010010001000100011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101111011011101110111011101110111011101011100100010000100100010001000100110110111011101110111011101110111011101110111011101,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100001100110011001100110011001100110100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010001000100010001010100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101100110010101100110011110001000100110011010101010101001100110011001100110011000100010001000100010001000011101110111011101110111011101110111011101111000100010001000100010011001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101111111111111111111111111111111111111111111111101111111111101111111111111111111111111111111111111111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011111101010000010010001000010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100000100010000100100010001000100101110011011101110111011101110111011101110111011101,
	2400'b001100110011001100110011001100110011010001000100010001000011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110011001101000100010001000011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001010101010101010101010101010110011001100110011001100110011101110110011101110110011001100110011001111000100110011010101010101011101110111010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001101110111011101110111101110111011101110111011011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111101111111111111111111111101111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110111111111110111011111110010100010001001000010010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100100010001000100010001000100100101011001100110011001100110011001100110011001100,
	2400'b001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101000100010001000100010001000011010000110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010110011001100101010101010101010101010101010101010101010101100110011001100110011001100110011101110111011101110111011101111000100010011001101010101010101010101010100110011000011101111000100110011001101010101010101110111011101110111011101110111011101110101011101110111011101110111011101110111011101110111100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110011000010001001000100010100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111110111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101100110010001000100010001000100011101011001100110011001100110011001100110011001100,
	2400'b001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010001000100010001000100010001000100010001000100010001000100010001000101010001000101010101000101010101010101010101010101010101010101010101000100010001000100010001000100010001000101010101010101010101010101010101010101010001000100010001000100010001000101010101010101010101010101010101000100010001000100010001000101010101010101011001100110011001110110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101111000101010111011101111001100101110111011101010011010101010101010101010101011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011011101110111011101110111011100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011100110011011101110111011101110111001100110011001101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101101111011101110111111101110111011111111111011101110111011101110111011101110111011101101110011001101111011101110111111111111111111111111111111101110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111011111110111011101110111011101110111011101110111011101110100000010001001000100010100011111111111111111111111111111111111111111110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110101000001000100100010001000100011100111011101110111011101110111011101110111011101,
	2400'b010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010001000100010001000101010101010101010101010101010101000100010101010101010101010101010101010101010101010100010001000100010001000100010001010101010101100110011001100110011001010101010101010101010101010101010101010101011001010101011001100110010101010101010101000101010101010101010101100110011001110111011101100111011101100110011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011110011010101110111011101111001100101110111011101110111011101110111011101110111011101110111100101110111100110011001100110011001100110011001100110011001011110011001100110011001100110111011101110111011101110011001100110011001100110011001100110011001100110011001100110010111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110111001101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101111111011101110111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101111111111111111111011101111111011101110111011101110111011101101110011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011110111011111111111111101111111011101110111011101110100100100001001000100001011111101111111111111111111111101110111111111110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110101100010001000100010001000100010100111101110111011101110111011101110111011101110,
	2400'b010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010001000100010001000100010001010101011001100110011001100110010101010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101100111011101110111011101110111011110001000100010001000100110011001100110011001100110011001100110001000100001111000101010111011101111001100110011001100110011001100110011001100110010111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011100110111011100110111011101110111011101110111011101110111011101110011001100101110111100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101111111111101110111011111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101111111111111110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111110111011101110110011001110111011101110111011101110111011101110111011101110101000100001001000100001010111011110111011101110111011001100110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110101110010001000100010001000100010011111101110111011101110111011101110111011101110,
	2400'b010001000100010001000100010001000100010001010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010100010001000100010001000101010001010101010101010110011001100110011001010110010101010101010101010101010101010101010101010101010101000100010001000100010001000100010101100110011101100110011101110111011101110110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101111000100010011001100110101010101010101010101010101010101010101010101010101010101010011001101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001011101010111011101111001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111101110111011111111111011101110111011101110111011101110111011111110111011111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110010111101111011101101110111001011101110111011101110101010101010101010101010101010101010101011100100100001001000100001010011001100110011001100101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001110110111001011101111001100110011001100110011001101110011011101110111011101110111011100110011011101110111011101110111011101110111101110111011101110111011101110111011101101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110101110010001000100010001000100010011011101110111011101110111011101110111011101110,
	2400'b010001000100010001000100010001000100010101010101010101010101010101010100010001000100010001000101010001010101010101010100010001010100010001010101010001000100010001000100010001000100010001010101010101000100010101010101010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010110011001100101010101010101010101010101010101010101011001100111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100110011010101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111101101111011101101110111011100101110101001100010011011110010111011101111001100110011001101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011111110111011111111111111111111111111111111111111111111111111111111111111111110111111101110111011101110111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011101010011011110011001100110011011100110011001011101110111011101110111011101110111011101110111011101000110001001000100001010011001110110111011101110110111011110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111101110010101010101010101010101010101010101010101010101010101010101010101010101110111010101010101011101110111011101110111011101110111011110010111011110011001100110011001011110011001100110011001100110011001100110011011110110111011101111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110000010001000010010001000100010010111011110111011101110111011101110111011101110,
	2400'b010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010011001100110011001100010001001101010101010101010101011110011001100110010111011101110111011110010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110011001101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110110111001010100010001000011110001000100110011001101111001100110011011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111101111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101110011001101110111101110111011101111111011101110111011101110111011101110111011101110111011101110110101000001000100100001001111001111111111111111111011101101110111101110111011101110110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110010111100101110111011101110111011101010101011101110111011100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101111011101101110111011101110111100110011001100110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110010010011001000100010001000100010010111011110111011101110111011101110111011101110,
	2400'b010001000100010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101100110011001010110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100101011001100110011001100110011001100111011101110111011101110111100010001000011110000111011110000111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010011010101010101010101010101011101110111011101110111011110011001100110011001100110011001011110011001100101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011011100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110110110111001100010001000100010001001100110011010110011011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100001000100010001001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110110111011110111011101110110111011101110111011101110111011100101010011010101010101010101010101010101010101010101010101011101010111011101110111011101110101010101010101001100110011001101010101010101010101010101010101010101010101010101010111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010111010101110101011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001011101110010011001000100010001000100010010010111101110111011101110111011101110111011101,
	2400'b010101010101010101010101010101010101010101010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101011001100110011001100110011001010101010101010101010101100110011101110111011110001000100010001000100010001000100010001000100010001000100001110111011101110111011110001000100010001000100010001000100010001000100110101010101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100101110111011101110111011101111001011110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110110111011101110111011101110111011101110010111001100110001000100010001001100110101011110011001100110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101110001001000100001001010101111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101101110111011101110011001100110011001100110011001100110011001100110011011101110111011101110010111011101110111010101010101011101010101010101110111010101110101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110101010101010010100001000100010001000100010001110101100110011001100110011001100110011001100,
	2400'b010101010101011001100110011001100110011001100110011001100110011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001110111011101111000100010001000100010001001100010001000100010001000100010001000100001110111011101111000100010001000100010001001100110001001100110101010101010101011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011100110111011101110111011100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011010101010101011110011001100110111011101110111001011101010011000100010011010110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111110000010001000100001001010011111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101101110111011110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100101110111011101110111011101110101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101001000100010001000100010001010001100101110111011101110111011101110111011,
	2400'b011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011010101010101010101010101010101010101010101010101011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011011100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101001110111011101110111100010001000100110011010101010011001101010101010101010111100110111011110111011101110111011101110111011101110111011101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111111101100101110111101111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110010010001000100001001010001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110110110111000100010101100110111011101110111011101110111011101110111011101110111011101110111001100101111001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100101110111011101110111011101110111011101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110010110001000100010001000100001001001111010101010101010101010101010101010101010,
	2400'b011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110110111011101110111011101110011001100110011001100110010111011100101110111011101110111011101110111011101110111011101110111100010001001101011001100110011011101110011011101110111011110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111110111011101111111011111111111111101111111010100111011110001001100110011001100110011011101110111100101110111011110111111111111111111111111111111111111111111111111011111111111011111110111011101110111011101111111011111111111011101110111011101110111011101110111111101111111111101111111011101110111111111111111111111111111111111111111111111111111111111111111110110010001000100001001001111110111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110101001110110011001100110100010111101110011011101110111001100110111001100110010111001100110011000011110001000101010111100110011001101110111011100110111001100101111001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111100110010111011101110111011101110111011101111001100110011001100110011001100110011001011101110111010101010101001100110011001100110011001100110011001100110011001100110000110001000100010001000010010001001101010101010101010100110011001100110011001,
	2400'b011001110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110010111011101110111011101110111011101110111011101010011000100010001000100110011001100110011001100110101010101010011010101010101011110011001100110011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111011101110111011111111111011101110111111111111111010010110011001111000101110111010100110001000100010001000100110101011110111101110111011101110111011101110111111111110111111101110111011111110111011111111111111111110111011101110111011101110111011101110111011101110111011101110111011111111111011101111111111101111111111111111111111111111111111111111111111101110111110110011001000100001001001101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111110111011101110111011101110111011101011011101100110011001100110011001111001100110101010101010011001100110011000100001110110010101010101010101010110011010001001100110101010101010101010101010000111011101110111011110101011110011001100110011001100110010111011101110111011101110111011101110111011101110111011110011001011101110111011101110111011101110111011101110111100110011001100110011001100110011001011101111001100110010111011101110101010101010101010101010101010101010101010101010100111001000100010001000010010001001011010101010101010101010101010101010101010,
	2400'b011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001001100110011001100110011001100110011001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111001100110011011101110011001100101110111011110011001100110011001100101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101001100110011010101010011010101010101011101111001100110011001100110011001100110011011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111010111000011101111000101010111100101110101010101110111011110011011110111111111111111111111111111111111110111011111111111111101110111011111111111011101111111111101110111011101111111011101110111011101110111011101110111011101110111011101111111011111111111111101111111111111111111111111111111111111111111111111110111111000011000100100001001001011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111101110111011101110111011101110111011101110111011101110111011001000011001100110011001100110010101010110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101100110011001100110010101010101010101010101010101111000101010111010101010011000100010011001100110001000100010001000100010001000100010011100110111011100101110111011101110111011101110111011101110111011101110111011101110111011101010001000100010011001101111001100101110111011101110111011101110111011101110111011101010101000001100100010000100010001001001001011110011001100110011001100110011001100,
	2400'b011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100110011001100110011010110011001010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111001100110111011100110011001100101110111100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010011001100110011000100010001000100010011001100110011001101010101010101110111100101111001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101111111011101111111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011011110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011111110111111111111111111101111111111101110111111010100001000100001000101001101111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010010111011001100110011001100101011001010110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011101110110011001010101010101010101010101010101010101010101010101010101011001111001101110111011101110111011101110111011101110101010101010011001100010001000100010001000011001010110011001110111100010111100101110111011101110111011101110111011101110111011101110111001001100100010000100010010001000111011110011001100110011001100110011001100,
	2400'b100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011010111011011010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100101110111010100110011001100110011001100110011001100110011001100110011001101010101011101110111011101111001100110011001100110111011101110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111100101001000100001000101001100111111111111111111111111111011111111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100101010001000011101110110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011101110111011101110111011101110110011001100110010101010101011001100101010101010101010101010101011001111000100010001000100010001001101010101010101110111011101110101001010000100001000100100010001000111001101010101010101010101010101010101010,
	2400'b100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101001110111011011101010111010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001011110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110011001100110011001100110011001100110011011101110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100101110111011101110111010101010101001100110011001100010001000100010011001100110011001100110011010100110101010101110111010101110111011101111001011110010111011101110111100101110111011110011001100110011001101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000010001000100111100111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101101110010111010100110011001011101100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100101010101010101010101010101010101010101010101010100010001010101010101010101010101010101010101100110011001100110011001110111100010011001101010101001010000100010001000010001000100100111100110011001100110011001100110101010,
	2400'b101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010110111011011101010111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101010101010100110011001100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100010011001100110101011101110111100110011001100110011001100110011001100110011011101110111011100110011001100110011001100110011011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100111001000010001000100101011111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001011101110111010101010010111011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000101010101010101010101010101010101010101010101010101010101010101010101100110011101110110010000100001000100010001000100100110100110011001100110011001100110011001,
	2400'b101110111011101110101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111001101010111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110010111100110011001011101110111011101110111011101110111011101110101010100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011011110011001100110011001011101010101011101111001100110010111011101110111010100110011001100110011010101010101010101010101011101110111011101110111011101111001100110011001100110011001101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111010111000100010001000100101001111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111101101110111011101110111011101110111001011101110101010101010101010100110011001100001110111011101100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010001000100010101010101010101010101010101010101010101010101010101010101010001000101010101010100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001000100010001000100100101011101111000100010001000100010001000,
	2400'b110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001101010111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101111001100110011001100110011001100110011001100110011001100110011001100110010111011101111001100101110111011101110111100101110111011101110111011101110111010100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010101110111100110010101001100110011001101010101011101110011001100110011001100110001000100010001000100010011001100110011001100110101010101010101011101110111011101110111100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110011001100101110111011101110101010101010100111000100010001000100101000110111011101110111001100101110111011101110111011101110111011101110111011101111001100110011001100110111001100110011001100101110101010100110011001100110011000100001110111011101110111011101110111011101110111011001100110011001100110010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000101010101010101010101010101010101010101010001000101010101010100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100010000100100001000100100100011001100110011001100110011001100110,
	2400'b110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011100110010111011101110111011101110111011101110111011101110111011110011001100110010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101111001100110011001100110011001011101110111100110010111011101110101001100110011000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100110011001100110001000100010001000100010011001100110001000100010001000100110011000100010001000100010001000100110011001100110011001100010011001101010111011101110111011110011001100101111001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110111011101110111011101110011001100110011001100101110111011101110101010101010101010101010101010101010101010101010101010101010100111000100010001000100010110101010101010101010011001101010011010101010101010101010101010101010101010101010101010101110111010101110111011101110111011101010101010101010101010101010011001100010001000100010001000100110011001100110001000100010000111011101110111011101110111011101100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010100010000100010000100100001000100100011010101010101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011011101110111011101110111011101110111101110110111011101110111011101110111001100101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111010101010011001100110001000100010001000100010001000100010001000100001111000100010000111011101110111011101110111011110001000011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010011010101110101000100010001000100010001001100110011001100110011010101010011010101010101010101111001100110011011101110111011101110111011101110111011101110111001100110011001100110011001100110010111011101111001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111001001000010001000100010100100110011010101010101010101010101011101010101010101010101010101010101010101010101010101010101010100110011001100110101010101010101010101010101010101010101010101010011001101010011001100110011001100110011001100110011001101010101010101010011001100110011001100110011000100010001000100001110111011101110111011101100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101000100010001000101010000100001000100010001000100010011010101010101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110111011101110111001101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111001101110111011100110111011101110111011101110111011110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001011101110111011101110111011101110111010101010101011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111100110011001100110011001100110011001100110011001100101110111010101010011001100110011001100110011001100110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100001110111100010001000100010001001101110111000011101110111100010000111011101110111100010001000100110011001100110011001101010111011101110111011101111001100110011001100110011001011101110101010101010111011101111001100110010111011101111001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111010001000010001000100010100101010111011110011001100110011001011101110111011101110111011101110111011101110111011101110111011101010011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110101010100110101010101010101010101010101010100110011000100010001000100010000111011101110111011101110110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100100001000100100011010101010101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110111001101110111011101110111011101110111011101110111011100110011001101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110011011100110111011101110111011101110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110010111011101111001100110011001100110011001100110010111011101010101010101111001100110011001100110010111011101110111011101110111011101110111010100110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111010101010101010101010111011101010101001100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100110011000100010000111011101110111011101110111011101110111100010001000100010011001101010101001100110011001100110101010101010101010101010101001100110011001100110011001101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010001100010001000100010011101111001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110101001100110011001100110001000100010011001100110101010101010101010101010101010101010101010101010101010100110011010101010101010101110111010101010111011101110111010101110111011101010101010100110011001100110011001100010001000100010000111011101110111011101110111011101110111011101100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001110111011001010101010101010101010101010100010001000100010001000100010001000100010101000100010000100010000100010001000100010011010101010101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111001100110011001011101110111011101110111011101110101010101010101001100110011001100110011010101010011010100110011001100110011001100110011001101011001100110011001100110011001100101110111011101110111011110011001010100110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101111001100101110111011101010011000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101111000100010001000011110001000100010001000100110011001100110101010100110001000100010001000100010001001100110011001100110101011101110101010101010101010101010101010101010101010101010101010101010101010101010111011101110101010101110111011101010101010001100010001000100010010100111001100110011001011101110111011101110111010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011000100010011001100110011001100110011001100110011000100010001000100010011001100110011010101010101010101010111011101110111011101110101010100110011001100110011001101010011001100110001000100010001000100010001000100010011001100110001000011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011001100110010101010101010100110001000100010001000100010010010101010101010101010101010101100110,
	2400'b101110111011110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011001011101110101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001101010111100110011001100110011001100110011001100110011001100110011001010101010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111001100110011001100110011001100110011001100110111001100110011001100110011001100110011001100101111001100110011001100110011001011101010011000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010011001100110011000100010001000100010001000100010001000100010011010100110011001100110011001100110011001100110011001100110011000100110011001100110011001101010101010101010101010101010011001001100010001000100010010011110101010101010101010101010101001100110011001100110011001100110011001100110001000100010011001100110011010101010101010101010101010101010101010100110000111011101110111011110001000100010001000100010001000011110001000100010001000100010001000100010001000100010001001101010101010101010011001100110011001100110011001101010101001100110011001100001110111011101111000100110101001100010001000100010001000100010001000100110011001100110011000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101111000100010001000100110011001100110011001100110011001100110011001100001110111011001100110011000110010000100010001000100010010010101100110011001100110011101110111,
	2400'b101110111011101110111011101110111100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011010101111001100110011001100110011001100110011001100110011001100110011001010101010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111001100110011011101110011001100110011001100110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001101110111011110111011011101110011001011101110111011101110111011101110111011101010101010101010101010101110111010100110001000100010001000011101110111011101110111011101110111011001100110011001100110011001100110011001100110011110001000100010001000011101110110011001100110011001100111011101110111011101110111011101110111011101111000100110011001100010001000100010001000100010001010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010000111001100010001000100010001011110011001100110011000100001110111011001110111011101100110011101110110011001100110011001100111011101110111100010001000100010000111011101110111011101110110011001100101010101010101010101100110011001100110011101111000100010001000011101110111011101110110011001100111011110001000100010011001100110011001100110011010101010101001100110000111011101100110011001100110011001110111011101110111011101110111100010001000100110101010101010101010101010101010101010101010101010111011101110101010101010011001100110001000100010001000100010001000100010001000100010001001101110111011101010101001100110011000100010001000011101110111011101110111011101000010000100010001000100010010011010001000100010001000100010001001,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101111001100110011001100110011001100110011001011101110111011101110111011101110101010101110111011101110101010101010101010100110011001100110011001100110011001101010101010101010101001100110011001100110011001100110011001100110011001100110101011110011001100110011001100110011001100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110111011101110111011100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110111011110111011101110111011101101110111011101110111011101110111011101110111011101110111011110111011101101110111011100110011001100110011001011101110111011101110101010100110000111011001100110011001100110011001100111011110001000011101110111011101100110011001100110011001100110011001100110011101110111011101110111011101110111100010011001100010001000100010001000100010001000100001110111100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110010000010001000100010001010110011001100110000111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101011001100110011001110111011101110111011101110111011101100110011001100110011001100111011101111000100010011001100110101010101010101001100001110111011001100110011001100110011001100110011001100110011001100110011001110111011110001000100110011001100110011010101010101010101010101010101010101001101010101010101010011001100110011001100110011000100010001001100110011010101110111010101010101010101010011001100110011000100010001000100010001000100001010010000100100001000100010001011110011001100110011000100010001000,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011001101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101001100110011001100110011001100110011000100010001000100110011001100110011010101010111011101110111010101010111011101111001100110011001100110011001100110011001100110011001100110011001100110011001010101010111100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011011101111011101110111011101110111011011101110111011101110111011101110111011101110111011110111011101110111011101110110111011101110111011101110111011101110111011101110010111001011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011110001000011101110111011101110111100010001000100010001000100010001000100010001000011101110111011101110111011001100110010000010001000100010001010010001000100001110110011001100110011001100101011001100101011001100110011001100101011001100101010101010101011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101011001100111011101110111011001100110011001100101010101010101010101010101010101010110011001100111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011110001000100010001000100001111000100010001000100110011001100110011001100110011001100110011001101010101011101110111010101010101010101010011001100110011001100110011001100110011000100001100010000100010001000100010001010110011000100010000111011101110111,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110011001100110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101111001100110011001100101111001011101110111011101110111011101110111011101110111010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110101010101111001100110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001010101011001100110011001100110011011101110111101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011111110111011011101110111011101110111011101110111011101110011001100110011001011100110000111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001100110011101110111011101110111011101110111011101110111100010000111011101110111011101110111011101110111011101110111011110001000100010001000100010001000011101110111011101111000011101100110011001100110010000010001000100010001001101111000011101110110011001010110011001100101010101010101010101100110011001100101011001010101010101010101010101010101010101010101010101010110011001100110011001010101010101010101010101010101010101010101010101100111011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010101010101010101010101010101010101010101011001010101011001100110011001100110011001100110011001100110011001100110011101110111011101111000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010001000100010001000100001100010000100010001000100010001001101110111011101110111011101100110,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011100110111011100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110111001100110011001100110011001100110011001100110010111100110011001100110011001011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111100110011011101110111011101110111011101110111011101110111011101110111011101110011001100110111011101110011001100110011001100110011001100110111001010101011001100110011001100110111011101110111101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110110111011101110111011101110111011101110111011101110111011100110011001100101110101001100010000111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101100110011001100110010000010001000100010001001101100111011001100110011001100101010101010101010101010101010101010101011001100110010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010101010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001110110011001110111011101110111011101110111011101110111011101110111011001110111011001110111011101110111011101110111011101100011000100010001000100010001001101100110011001100110011001100110,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100101110111011110011001100110011001100110111011100110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001011101111001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101010101001100110011001100110011001100110011001101010101011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011110011001100110111011101110111011101110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001010101011001100110011001101110111011101110111101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011011101111011011101110111011101110111011101110111011101110111011110111011101101110111011101110111011101110111011101110111011101110111011101110111011110111011101110110111011101110111011101110111011101110111011101110111011101110011001011101110111010100110011000011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110110011001100110011001100110011001100101010100100001000100010001001001100110011001100110011001100101010101010101010101010101010101010101010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010101010101000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100011000100010001000100010001001001010101011001100110011001100110,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011100110011001011101110101010101010101001100110011001100110011001101010101001100110011001100110011000100010001000100110011001101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110101011101110111010101010101001101010101010101010101010101110111011101110111011101110111011101110111011101110111010101010101001100110001000100010001000100010001000100010001000100110011010101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011010101010111011110011001100110011001011101011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001010101011001100110011011101110111011101110111011110111011011110111011011101110111011101110111011101110111011101110111011101110111101110111011101110111011101101110111011101110111101110111011101110111011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011110111011101110111011011101110111011101110111011101110111011100110111011101110111001100110011001011101010011001100010000111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110110011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010100100001000100010001001001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101010100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000101010101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001010101011001010101010101010101010101010101010101010011000100010001000100010001001001010101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101010011000011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011110001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011000100110101010101010101010101110111011110011001100110011001100110011001011101110111011101010101001100010001000100010001000100010001000100110011001100110011001101010101010101010111011101110111011101110111011101110101010101010111011101110111011101010101010101010101010101010101000100010001000100010011001100110001000100010011001101010111011110011001100110011001011101011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001010101011001100110011011101110111011101110111011110111011101110111011101110111011011101110111011110111011101110111011101110111011101110111011101110111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011101110110111011101110111011101110111011101110111011101110111001100110011001011101110101001100110011001100010001000100001110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010100100001000100010001001001010110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001010101010101000100010001000100010101010101010101010101010101010101010101100110011001010101010101010101010101010101010101010101010101010101010101010011000100010001000100100001001001000101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111010100110000111011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001110111011101110111011101110111011110001000100010001000100010001000100010001000100001110111100010101010101010101011110011001101110111101110111011101101110111011101110011001100101110111010100110001000100010001000100010011001101010111011101010101010101010101010101010101010101010101010101110111011101110111011101110111011101010101010101010101010100110011001100110000111011110001000100010011001100110011000100010011001101110111011110011001100110011001011101011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001011101111001101110111011101110111011101110111101110111011101110111011101110111011101110111011101101111011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111011101110111011101101110111011101110111011101110111011101110111001100110011001100110011001010101010011001100110101010101010101001100110000111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010100100001000100010001000101010110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101000101010101010101010101010100010101000100010101000100010001010100010001000100010001000100010001000100010001000100010001000100010001000101010101000101010001000101010101010100010001010101010101010101010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101100110010101010101010101010101010101010101010101010101010101010011000100010001000100100001001001000101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110101001011101100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000011101100110100010011001101010101010101110111100110111011110111011011101110111011100110011001100101110111010100110001000100010001001100110011001100110101010101010101011101110111011101110101010101010101010101010101010101010111011101110111011101110111010101010011001100110001000100001110111011101111000100010011001100110011000100010011010101110111011110011001100110011001011101011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001011101111001101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011101110111011101101110111011101110111011100110011001100110011001100110010111011101010101010101110111011101110101010100110011000011101110111011101110111011001100110011001100110011001100110011001100110011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010100100001000100010001000101000110010101100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010001010100010001000100010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010110010101010101010101010101010101010101010101010101010101010011001000010010001000010001001001000100010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110101001011101100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100111011101110111011110001000100010001000100010001000100010011001100010001000100001100110011110011001100110011001101010101011110011001101110111001100110011001100101110111011101110101010101010011001100110011001100110011001101010101011101010101010101010111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010011001100110011000100010001000100010011001100110011001100110011010101110111100110011001100110011001011101011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011011101110011001011101110111011101010101010101010101010101010101010101010011001100110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001010101010101010101010101010101010100110001000100010001000101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001010100010001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010001010100010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010100010101010101010101010101010101010101010101010100000100010010000100010001000101000101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111010100001110110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001110111011101111000100010001000100010011001100110011001100110011000100001100110100010101010101010101010101010101011101110111011101110111011101110111011101010101010101010101010101010011001100110011001100110011010101110111011101010101010101010101010101010101011101110111011101110111011101110101010101010101010101010101010101010101001100110011001101010011000100010001000100010011001100110011001100110011010101110111100110011001100110011001011101011001101110111011101110111011101110111011101110111011101110111011101110111011101110111001011101111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011101110111011101110111011101110111011101101110111101110111011101101111011011101110011001011101110111011101110111010101010101010101010011001100110011001100110011000100010001000011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001100101010101010101010101010101010100110001000100010001000101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010100001000010001000100010001000100110101010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110011011101110111001100110011001100110011001100110011001100110011001011101010000111011001100101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001110111011101111000100010001000100010011001100110011001100110011001100001100110100010101011110010111011110011001011101110101010101010101010101010101010101010101010101010101001100110011001100110011001100110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101110111011101010101010101010011000100010001000100010011001100110011001100110011010101111001100110011001100110011011100101111001101110111011101110111011101110111011110110111011101110111011101110111011101110111011011101111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110010111011101010101010101010101010101010101010101010101001100110011000100010001000100001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010100110001000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010100001000010001000100010010000100110100010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110011011100110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001011101010011001100001110111011001100110010101010101010101010101010101010101010101010110011001100110011001100111011101111000100010001000100010001001100110011001100110011001100001100110011110001001100110011001100110101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101001101010101010101010101010100110011001100010001000100010011001100110011001100110011010110011001100110111011101110111011101101111001110111011101110111011101110111011101110111011101110111011101110111011101110110111011011110011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110010111011101010101010101010101010101010101010101010101001100110011010101010101010101010001000011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101000001000100010001000100110101010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010001010100010001010101010101010100001000010001001000100010000100110100010101010101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111001101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100101110111011101010011000011101110110010101100101010101010101010101010101011001100110011001100111011101111000100010001000100010001001100110011001100110011001100001100110011110001000100010000111011101111000100010011001100110011010101010011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010100110011001100110001000100010001000100010001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001100110101011110011011101110111101110111011101101110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011011011110011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011101110111011011101110111011101110111011101110011001100110011001100110011001100110011001100101110111011101110111011101110111011101010101010100110011010101010101010101010101010100110011001101010101010101010011001100010001000100010001000100010001000011101100110011001100110010101100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101000001000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010100001000010010001000100010000100110100010001000101010101010101,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110011001101110111011101110111001100110011011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110010111011101110111010100001110110011001100110011001010101010101100110011001100110011001100111011110001000100010001000100010001000100010011001100110011001100001100110011101111000100010001000100010000111011101110111100010001000100010001001100110011001100110011001100110011001100110011010101010101010101010101010101010011001100110011001100010001000100010001000100010011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010100110101010101010011001101010101011110011011101110111011110111011101101110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011011011110011011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101111111111101110111011101110111011101110111011101110111011101110111011011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110101010100110011001100010001000100010001000100010001000011110001000100010001000100010001000100001110111011101110111011001100111011101100110011101110111011101110110011001010101010101010101010101010101010101010101010101000001000100010001000100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010001010100001000010010001000100001000100110100010001000100010001000100,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111001101110111001100110011001100110011001100110011001100110010111011101010101010101010101010100001100110011001100110011001100110011001100110011001100110011001100111011110001000100010001000100010001000100010001000100010001001100001100110011001100111100010001000100110011001100010001000100010000111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010100110101011101010101010101010101011110011011101110111011101111011101101110011011101111011101101110111011101110111011110111011101101111011101110111011101110111011011011110011011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110010111011101110111010101010101010100110011001100010001000100010001000100001110111011101110111011101110111011101111000100010001000100010001000100010001000011101110111011001100110011001010101010101010101010101010101010101010101010101000010000100010001000100100101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100001000010001000100010001000100100100010001000100010001000100,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111010100010000111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100111011101111000100010001000100010001000100010001000100010001000100001100110011001110111011101100111011101110111100010001000100010001000100010001000100001110111011101110110011001100111011001100110011001100111011101110110011101110111011101110111011101110111011110001000100010001000100010001000100110011001100110011001101010101010101010101010101010101001100110101001100110101010101010101010101010111011110011011110111011101110111011101110110111011110111011101110110111011101110111011101110111011101111011101110111011011101110111001011110011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110111011101110111011101110111011101111111111111111111111111110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110010111011101010101001100110011000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110010101010101010101000010000100010001000100100101010101010101010101010101011001010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100001000010001000100010001000100100100010001000100010001000100,
	2400'b110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110101001100010000111011001100110010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001110111011110001000100010001000100010001000100010011010101010011001100110101010100001110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011110001000100010001001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101111001100110011011110111011101110111011101110110111011101111011101110111011101110111011011101110111011101110111011101110111011101110111001011101111001101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101111011101111111111111111111111111111111111101111111011111111111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100101110111010101010101010101010101010101010101010101010011001100110011000100010000111011101110111011101100110011001100110011001100110011001100110011001100110011001010101010101010101010101010010000100010001000100100100010101010101010101010101010101010101010101010101010001000100010001010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101010101001100010000111011101100110011001010101010101010110011001100110011001100110011001100110011001100110011001111000100110011000011101110110011110011010101010101010101110111011101010011001100110011001100001110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011110001001101010101011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010111010101010101010101010101010101010101011101110111011101111001100110011011101111011101101110111011101110111011101110111011101110111011101110111011101110111011100110111011101110011001100110011001100110011011101110111011101111011101110111011101110111011101110111011101110111011101101111011101101111011101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110011011100110011001100110111001100110011001100110011001100110011001100101110111011101010101010100110011001100010001000100001110111011101110111011101110111011101100110011001100110011001010101010101010101010101010010000100010001000100010100010101010101010001000101010001010101010101000100010001000100010001010101010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111010100110011000100010000111011101110111011001100110011001100110011001100110011001100111100010011001100110000111011101111000100010001000100010011001100110011001100110011001101010101010100110011001100110001000011101110110011001100110011001100101011001100110011001100110011001100110011001100110011001100111100010001000100010011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010011001100110101010101010101010101010101010101010101011101110111100110011011100101110111011101110111011101110111011101110111011101110111100110111011101110111011101110011001100110011001100110111011101110111011101110111101101110111011110111011101110110111011110110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011101111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111101110110111101110111011101110111011101101110111011100110011001100101110111011101110111011101110111011101111001011101110111011101110101010101010101010101010101010101010101001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100011000100010001000100010100011001010101010101010101010101010101010001010101010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011010001000100010101010101010101010100010001010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101010101010100110011000100001110111011101100110011001100111100010001001100110011000100110001000100110011000100010001001100110011001100110011001100110011001100110101010101010101010101010011001100110000111011101100110011001100101010101010101010101100110011001100110011101110111011101100110011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100110011000100110011001100110011001101010101010101110111011101010101010100110011001100110011001100110011001100110101011110011011101110111011101110010111011101110111100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101101110111011100110011001100101110111011101110111011101110111011101110111011101110111011101010101010100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110100000100010001000100010100100001110111011101110111011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010001000100010001000100010001010101010101010101010001000100010001000100010001000100010001000100010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100001100110011010001000101010101000101010101010100010001010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111010101010101010100110011000100010001001100110001000100010001000100010011000100110101010101010101001100110011001100010001000100010001000100010001001100110011010101010101010100110011000011101110110011001100110011001100110011001100111100010001000100010001000100001110111011101100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111100010001000100110011001100110011001101010101010101010101001100010001000100010011000100010001001100110011001101110111100110010111011101110111011101010111011101110111011101111001101110111011101110111011101110111011101110111011101110111011101110011011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111101110111011101110110111011101110111011101110011001100110111011101110111011101110111011100110011001011101110101010101010101010101010101010100110011001101010101010101010101010101010101010100110001000100010000111011101110111011101110111011101110111011101110101000100010001000100010100100110011001100110001000100010000111011101110111011101110110011001100110011001100110011001100110011001010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010001000100010001000100010001000011001101000100010001000100010001000011001100110011001101000100010001010101010101000100010001000100010001000101010001000100010001000100001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101010101010100110011001100110011000100010011001100110011001101010101010101010101001100110001000100001110111011101110111011110001000100010001000100010001000100001110111011101110111011101110111011101110111011110001000100010001000100010001000011101110110011001100110011001100110010101010101010101100110011001100110011001100110011001100110011001100111011101110111011110001000100010001000100110001000100010001000100010001000100010001000100010001000100010001000100110101011101110111011101010101010101010101010101010101011101110111011110011001101110111011101110111011101110111001100110011001011110010111100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011011101110111001100110011001100110011001100110011001100110011011101110111101110111011101110110111011101110010111011101010101010101010101010101010101010101010101011101110111100110011001011101110111010101010011001100110001000100010001000100010001000100010000110000100010001000100010100100010001000100010001000100010001000011101111000100001110111011001100110011001100110011001100110011001100110011001100110011001010110010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010001000100010001000100010001000100010001000100010000110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111001100110011001100110001000100010001000100110011001100110011010100110011001100010001000011110000111011101110111011101111000100010001000100010001001100110011001100110011001100110001000100010001000100010001000100010001000100010000111011101110111011001100110011001010101010101010101010101100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011110001000100110011001100110011001100110101001100110011010101111001100101110111010101010111011101110111010100110011000100010011001100110101100110011001100110011001100101110111100110011001100110011011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111001100110011001100110011011101110111011101110111011110111011101101111011101110110111011100110010111011101110111011101110111100110011001101110111011101110111011101110011001100110011001011101110111011101010101010100110011001100110010111001000010001000100010011011110000111011101110111011101110111011101110111011101110111011001100110011001010101010101010101010101100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010001000100010001000101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101000100010001000100010001000100010001000100010001000011001100110011001100110011001100110100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101010101001011110001000100010001000100010001000100110011001100110011001100110011001100010001000100010000111011101110111100010001000100110011010101010101010101010101010101010101010100110011001100010001000100010001000100010001000100010001000100001110111011001100110011001010101010101010110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101100111011101111000100010001000100010001000100010001010101110111100101110011000100010001000100010001000100001110111011110001000100010111100110011001100110010111010101010101010101010111100110011001100110011001100110011001100110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011011110110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101101111011101110111011011101111011101110111011101110110111101101110111011100110011001100110111011101110111101110110111011101110111001100110011001100110011001100110010111011101110111011101110101010101010101000001000010001000100010011011110001000100010001000011101110111011101110111011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011010001000100010001000100001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100110011001100110011000100010001000100001110111100010001001100010011001100110011001100110011001100110011000100010001000100010011001100110011001101010101010101010111011101110111011101110111010101010101001100110011001100110011001100110011000100010001000011101110111011001100110011001100101010101010101011001100110011001100110011001100110011001100110011001100110011101110111011101110110011001100110011001100110011001100111011101110111011101110111011101111000100010001000100001110111011101110111011110001000100001110111011101110111100110111100110011001100110010101001100110011001100110101010101110111011101110111011101111001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011011110111011101110111011101110111011101111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110011001100110010111011101110111011101110111011101110111011101010101010100110011001100110011000001000010001000100010010011110001000100010001000011101110111011101110111011101111000011101110111011101110110011001100110011001100101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010000110100001100110100010001000100010001000100010001000100010001000100010001000100001000010001000100100001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111010101010101001100001110111100010001000100010001000100010001000100010011000100110011001100110011001100110011001100110011001100110011001101010101010101010101010101110111011101110111011101110111011101010101010100110011001100110001000100001110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101111000101010111100110011001100101110011001100110011001100010011001100110101011101110111010101010111011101110111011101110111100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011011110111011101110111011101110111011101111111111111111111111111110111111101110111011101110111011101110111011101110111011101110111011101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011110111011011101110111011101110111011101110111101110111011101110111011101110111011101110110111011101110011001100110011001100110011001100110010111011101110111011101110101010101010101010101010101010101010101010101010101001001100010001000100010010011110011001100110011001100110011001100110101010101010111011101110111011101010101001100110011000100010001000011101110111011101100110011001100101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101000101010101010101010101010110011001100110010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010001010101010001000100010000110011001100110011010001000100001101000100010000110100001100110011001100110011001101000100010001000100010001000100010001000100010001000011001000010001000100010001000100010100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110101001100110011001100110001001100110001000100110001000100010001000100010001000100010011001100110011001101010011001101010011001100110011001101010101010101010101011101110111011101110111011101110111011101010101010100110001000011101110111011101110111100010001000100010000111011101110110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010110011001100110010101010101010101100110010101100110010101010101010101100110011001100111011101110111011110001001101110101010101110111010100110011000100110011001100110001000100110011001101010101011101110111011101110111011101010111011101111001100110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011011101110111011101111011101110111011101110111011101110111011101110111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011110110111101110111011011101110111011101110111011101110011001011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011010000010001000100010010011110111011101111001100110011001100110111011101110111011101110111011100110011001011101110111011101010101010101010011001100110011001100110001000011101110111011001100110011001100110011001100110011001100101010101100101010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010101011001100110011001010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010100010001000100010001000100001100110011001100110011001101000100001101000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010001000100100100010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011100110011001100101110101010101010011001100110011001100010001000100010000111100001111000100010001001100110011001101010011010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111010101010011000100001110111011101110111100010001000100110001000100010000111011101100110011001100110011001100110011001100110010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011101110111011110001011101010000111100010101001011101110111011101110111100110011000100010011001100110011010101110111011101110111011101110111011110011001100110011001100110011011101110111011101110111011110111011101110111011101110111011011101110111011101110111011101110111101110111011101110111011101110111011101110111011111111111111111111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110010111011101110111011101111001100110011001100110011011101110111011101110111011101110111011101110111011101110111001100110011001100010100010001000100010010011111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100101110111011101110111010101010101010101010011001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000010001000100010001001000100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110011001100101110111010101010011001100110001000100010001000100010001000100010001000100010011001100110011001100110011010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111010101010011001100010001000100010001000100010011001100110011001100110000111011101110110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011110011010101001110110011001110111011001100110011001100110011110001001100110001000100010011010101010101011101110111011101111001100110011001100110011001100110011001100110111011101110111011101110111101110111011011101110111011100110011001100110011001100110011001101110111011110111011101110111011101110111011101110111011101111111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001011101110101010101010101010101110111011110011001100101110111011101110111011110011001100110011001101110111001100110011001100110011001100110011001100110011001100110011001100010100010001000100010010011011001100110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100101110111011101110101001100110001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011000100010001000011101110111011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100101010101010101010101010100010001000100010001000100010001000100010001000100001100110011001100110011001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100001100110011010001000011001000010001000100010001000100100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111001100101110111011101010101010100110011000100010001000100010001000100010001000100010001000100010001000100110011001101010101010101010101010101010101010101110111010101110111011101110111100110011001100101110111011101010101001100010001000100110101010101010111010101010101010101010011001100010000111011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001111000100101100110011001100110011001100101010101100110011001100111100001110110011110001001100110101010101010101010101010101011101110111011101110111011101110111100110011011101110111011101110111011101110111001101110111011100110010111011110010111011101110111100110011011101110111011101110111011110111011101110111011101110111111111111111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110110111011101110111011101110111011101110111011100110011001100110010111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001011101110111011101110111011101110111100011100010001000100010001011011001100110111011101110111011101110011001100110011001100110011001011101110111010101010111011101110111011110011001100110011001100110011001100101110111011101010101010101010101001100010001000100010000111011110001000100010001000100010001001100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001010101010101010101010101010101010101000100010101000100010101000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010000110011010001000011001000010001000100010001000100100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100101110101010101010011001100110001000100010001000011101110111100010000111100010001001101010011010101010101010101010101010101010111011101110111011101110111011101111001100110011001100101110101010100110011010101010101010101110111011101110111011110010111011101110101001100110000111011101110110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100101011001100110010101010101010101010101010101010110011001100110011001111000100110011000100010000111011101111000100110011010100110011001100110011010101110111100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101111001101110111011101110111011101110111011101111011101110111111111111111111111110111011101110111011101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011100110011001100110011001100110011011101110111011101110111011101110111011100110111001100110011001100110011001100110011001101100000010001000100010001011011011101110111011101110111001100110011001100101110111011101110101010101010101010101010101010101010101010101010101010101010101011101111001011101111001100110011001100110011001011101110101010101010011000100010001000100010000111011101110111011101110111011101110111011101110111100010001000100010001000011101110111011101100110011101110111011101110111011101110111011001100110011001100110011001100101011001100101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010000110100010000110011001100110011001100110011001100110100010001000100010001000100010001000100010001000011001000010001000100100001001000100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100101110101000100010001000011110000111011101111000011101111000100010001001100110101010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110010111011101110111010101010101010101010111011101110111011101111001100110011001011101110111011101010101001100001110110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100111011101110110011001100110011001100110011101111000100010011000100010001000100010011010101110111100110011001101110111011100110011001100110010111011101110111011101110111011101110111100110111011101111011101110111011101110111011101111111111111111111111111110111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101100100100001000100010001011011101110111011101101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001011101010101010101010101010101010101010101111001100110011001101110111011101110011001100101110101010100110011000100010001000100010001000100010001000011101110111011101110111011101110111011101110110011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100101010101010101010101010110010101010110011001100101011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010100010001000100010001000011000100010001000100010001001000100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110010111010100110001000100010000111011110001000100001111000101010011000100110001000100110011010101010101010101010101011101110111011101110111011101110111011101110111011110011001100110111011100110010111011101010101010101010101010101110111011101110111011110011001100110011001100110010111011101010011000011101110110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100111100010001000011101111000100010001001100110011001101010111100110011001100110010111010101010101011101010101011101110111011101110111011110011001101111011101110111011101110111011101111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110111011101101110111011101110111011101110111011101110111001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001101101000100001001000010001010111011101110111011101110111011101110111011101110111011100110111001101110111011101110111011101110111011101110111011100110010111100101110111011101010101001100110101010101010111011110011001100110111011101110111011101110011001010100110011001100110001000100010001000011110000111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100111100010011001100110011001100110011000100001110111011101110111011001110111011101110111011101110110011001100110011001100110011001100110011001100111011101100110011001010101010101010101010101010100010001000100010001000011000100010001000100010001000100100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110010111010100110001000100010001000100010001000101010111010100110011001100110011001100110011010101010101010101010111011101110111011101111001100101111001011110011001100110011001101110111011101110111001100110010111011101110101010101010101010101010111011101110111011110011001100110011001100110010111011101110101010101010101011101110111011101110111011101110111010100110000110010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011101110111011101110111100010001000100010001000100010011001101010101010101010011001100110011010101010011001101010111100101110111011101110111011110011011101110111011110111011101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001101101100110001001000010001010011001101110011011101110011001100110011001100110011001100110011001100110011001100110011001011110011001100110011001100110011001100110011001100110010111011101010101010101010101010101010101010101110111011101110111011101110111010101010101010101010101001100110011001100110011001101010101010101010101010101010101010100110011001100010001000011101110111011101110111011101110111011101111000100010001000100010011001100110001000100010001000100010001000100010000111011101100101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100001100110011001100110011001100110100001100110011001101000011001000010001000100010001000100100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001011110010111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111101101110111011110110111011101110111011101110111011100110010111011101010101010100110011001100110011001100010011001100110101010101010101011101010101010101010101010101010111011101110111011101110111011101110111011101111001100110011001101110111011101110111011101110111001100101110111011101010101010101010101010101010101010101010111011101110111011101110101010100110011001100110011010101010101011101111001100110011001010011101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011101110111011110001000100001110111011110001000100010011001100010001000100010001001100110011001100110101011101110101010101010101010101010111011110011001101110111011110111011101110111011011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111100110011001100110011001100110011001101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111001100110011001100101100110001000100010001001110101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111101110111011101101110111001100110011001100110010111011101110101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101111001100110011001100110010111011110011001011101110111010101010011000100001110111100010001001100110101010101010111011101110101010101010011000011101110111011101110111011101110111011101110111100001110111011101110110011001100110011001010101010101010101010101000100010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000010001000100010001001000100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101111001011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011110111011101101110111011110110111011101110111011101110011001100101110111011101110111010100110011001100110011001100110101010101110101010101010011001100110011001100110101010101010101010101010101010101110111100110011001100110011001100110011011101110111011101110111011110110111011101110011001011101110101010101010101010101010101010101010101010100110011001100110011001100110011000100110011001100110011010101010101001100001110110010101010101010101010101010101010101010101010101010101010101010101010101011001100101011001100110011001100110011001110111011101110111011101110111100010001000011101110111011101111000100010001000100110011010101010101010101010101010101010101010101010111011110011011110111011101110111011101101110111011101110011001100110011001101110011011101110111001100110011011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111001100101110111011101110111100101110111011101110111100101101000001000100010001001010101101110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110011001100110011001100110011001100110010111011101110111011101110111011101110111010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110101010100110011000011101110110011001100110011001100110011001111000100010011001100110011000100001110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000011101110111011101100110010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000010010001000010001001000100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101111001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011110111011101110111011101110111011101101110111011101110111011101110011001100101110101010100110011001100110011010101010101010101010011001100110101010101010101010101010101010101010111010101010111011101110111011101110111100110011001100110111011101110111011110111011101110111011101110111011101110111011011101110111011101110111001100110011001100110011001100101110111011101110111011101010101010101010111011101110111011101010011000100001110111011001100110011001010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100111100001110111011101110111011101110111011101111000100010001000100110011010101010101010101010101010101010101010101110111100110111101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011100110010111011101110111011110011001100110011001100110001000001001000100001001010101101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001101110111011101110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110101010101010101010101010011001100110011001100110011000100010001000100010001000100010000111011101110111011101110111011101100111011101110110011001100110011101110111011110001000100010001001100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101100110011001100110011001100110010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000011001000100010001000100001001000100011010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100101111001011101110111100110011001011101111001011110011001100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011110111011101101111011101101110111101110110111011101110111011101110111011100110010111011101110101010101010101001100110011001100110101011101110111011101110111011101110111011101110111010101010111011101110111011101110111011110011001100110111011101110111011110111011101110111111111111111111111111111111101111111111101110111011101101110111011101110111001100110011001100110011001100110011001100110011001101110111011101110011001011101110101001100110000111011001100110010101010101010101010110010101100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111100010001001100110011001100110011001100110011010101010101010101110111100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011011101110010111011101110111011110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100010001001010101101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101010101010101010011001100110011001100110011000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101001100110011001100110011000100010001000100010001000100001110111011101110110011001110111011101110110011001100110011001010101010101010101010001000100010001000100010001000100010001000100010001000100001000100010000100100010001000100010010001000100010001000100,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110110111011101110111011101110111011100110011001011101110101010101010101010101010111011101110101010101010101010101010101010101010111011110011001100101110111100110011001100110011001100110011011101110111011101111011101110111011101111111111111111111011101111111111101110111011101110111011101101110111011101110011001100110010111011101110101010101110111100110011001100110011011100110011001011101110101001100001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101111000100010011001100110011001100110011001101010101001100110101010101010111011110011001100110111001100110011001100110111011101110111011101110111011101110111011101110111101101110111011101110111011100110010111011101010101010101110111011101110111011110011001100110011001100110011001100110011001100110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101111011101110111011101110111011101110111011101110110111011110110101100001000100010001001010011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101010101010101010101010101010011001100110011010101010111011101110111011101110111011101010111010101010101010101010111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101110111011101010101010100110011001100110011000100010001000011101110111011101110111011101100110011001100101010101010101010101010101010101010101010101010100001000010001000100100001001000100011011001100110011001100110,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110110111101110111011101110110111011101110111011101110011001100110011001100110011001011101110111011101110101010101010101010101110111011101110111011110011001011101111001100110011011101110111011101111011011110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011011101110111001100101110111010101010101001100110101010101010111011101110111100110011001100110010111011101010011000100001110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111100010001000100110011001100110011001100110011001100110011001100110101010101110111011110010111011101110111011101111001100110011001100110111011101110111011101110111011101110111001100110111001100110010111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110111011101110111011101110111011110110111101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111001110010001000100010001010001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100101110111011101110111100110011001100110011001100110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010011001100110011001100110011001100110011000100010001000100010001000100010001000100010000101001000010001000100010001001000100011011001110111011101110111,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101101110111011101110111011101110111011100110011001100110011001100101110111011101110111011101110111011101110111011101111001100110011001100110011001101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111001100101110111010101010011001100110011001100110011010101010101010101010101010101010101010101010011001100010000111011101100110011001100110011001100110011001100110011001100110011101110111011101110111011110001000100010001001100110011010101010011001100110011001100110011001100110101010101010101010101110111011101110111010101010101010101010101010101110111011110011001101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100101111001100110011001011101110111011110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001110010001000100010001001111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001011101110111100110011001100110011001100110011001100110011001100110010111011110011001100110010111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110001000100010001000100010011000100010000101001000100001000100010001000100100010011010000111011101110111,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101111011101111111111111111111111111110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011011101110111001100101110111010100110011001100010001000100010001000100010001000011110001000011110001000011101100110011001100110011001100110011001100110011001100110011001100111011101111000100010001000100010011001101010101010101010101010101010101001100110011001100110011001100110101010101010101010101010101010100110011001100110011001100110011001100110101011101110111011110011001100110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001011101010101010101010101010101110111011101110111011110011001100110011001100110011011101110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110110000010001000100001000101101100110111011101110111001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110001000100010001000100010001000100010000101001000010001000100010001000100100011011010001000100001110111,
	2400'b101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111001100110011001100110011001100110011011100110111011101110111011101110111011101110111101111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011100110010111011101010101010100110011001100010001000100010000111011101100110010101010101010101010101011001100110011101110111011101111000100010001000100010001000100110011001101010101010101010011001100110011000100010001000100010001001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001101010111100110011011101110011001100110011001100110011001100110011001100110011001100110011001100101110101010101010111011101110111100110011001100110011001100110011001101110011011101110111011101110111011101110111011101110111011101110111001011101110111011110011001101110111011101110111011101110110000010001000100001000101001011110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011011100110011001100110011001100110011001100110011001100110111001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101001100110011001100110011001100110001000100010001001100010001001100110011001100110011001101010101010101010101001100110011001100110011001100110101010101010101010101010101010101010101010100110011001100110011001100110000101001000010001000100010010001000100011011110001000100010000111,
	2400'b101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110101011101110111011101110111011101110111011110010111011101110111011101110111100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101111111111111111111111101110111011101110111011101110111011101110111011101110111011111111111011101110111111101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110011001011101110101010100110010111011101100110010101010101011001100111011110001000100010001000100010001000100010001000100010001001100110001000100010000111011101110111011101110111100010001000100010001000100010001001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010011001101010111100110011001100110011001100110010111011101110101010101010101010101110111011101111001011110011001100110011001100110011001011101110111011101110111011110011001100110111011101110111011101110111011110111011101110110111001010101010101001100110101010101111001101110111011101110110010010001000010001000100111010110010111011101110111011101110111011101110111011101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011110010111011101110111011101110111100110011001100110011001101111011101101110111001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110000101001000010001000100010001001000100011011110001000100010000111,
	2400'b100110011001100110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101111011011101110111011101110111011101110111011101110111011101110111101111111111111111111111111111111111111110111111111110111111111110111011101110111011101110111011101110111011101110111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111001100101110101001100001110111011101111000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101100110011001100111011101110111011101110111011101111000100010001000100010001000100010000111011101110111011101111000100010001000100010001000100010001000100010011010110011001100110010111011101010101001100110001000100010011001100110101010101110111011101110111011101110111010101010011001100110011001100110011001101010101011110011001101110111011101110111011101110111011100101110101010101010011001100110011001100110101010101111001100110110100010001000010001000100111010110011001100110011001100110011001100110010111011101110111011101110111100110011001100110011001100110011001100110011001100110111011101110011001100110010111011101110111011101010101010101010101010101010101010101110111011110011001100110011001011101110111011101111001100110011001100110011001100110011001100110011001100110011001011101110111011110011001011110011001100110011001100110011001100110011001100110011001011101110111011101110111011101111001100110011001100101110111011101110111011101110111010101010101010101010101010100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010000101001000100001000100100010001000100011011110001000100001110111,
	2400'b101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011110111011101111111111111111111111111111111011101110111011111111111111111111111011101111111111111110111011111111111111101110111111101110111011101110111111101110111011101110111011101110111111101110111011101110111011101110111011101110111011101110110111011101110111001100101110101001100010001000100001110111011101110111011101110111011101110111011101110111011001110110011001100110011001100110011001100110011001110111011101110111011101110111011110001000100010001000011101110111011110001000100010001000100010001000100010001000100010011011110111011100101110101010100110011001100010001000100010001000100010011010101010101001100110011000100010001000100010001000100010001000100010011001100110011001101010111100110111011101110111011100101110111010101010011001100110011001100110011001100110011001100110011010101010010010001000010001000100101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011110011001100110011001100110011001100110011001011101110111010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101001000100010001000100010001000100011011110001000100001110111,
	2400'b101010101010101010101010101010111011101110111011101110111011101110111010101010011001101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101110111011111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001011101010011001100010001000100010001000100010001000100010000111011101110110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100110101010101110111010100110011000100010001000100010001000011101111000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010001000100110101100110111011100110011001100110010111011101010101001100110011001100110011001100110011001100110011001100101110010000100010001000100101001110111001100110111011101110011001100110111011100110011001100101110111011110011001100110011001100110011001100110011001100110010111011101110111100110011001011101110111011101110111011110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111010101010101010101010101011101111001100110011001100110011001011101110111010101010101010101010101010101010101010101010101010101010101010101010101011101110101010101010111011101110111011101110111011101110111011101110111011101110101010101010100101001000100001000100100010001000100011011110011000100010001000,
	2400'b101010101010101010101010101010101010101010111011101110111010101010101000011101100110100010011001100110011001100110011001100110011001100110101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111011111111111111111111111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011100110011001100101110111010101010101010101010111011101110101000011101110110011001100110011001100101010101010110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111100010011010101010010111100010001000100010001000011110001000100010000111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101111000100010001000100010001010110010111010101011001100110011001100110010111010101010101010101010101010101010101010101010101001100110000011000100010001001000101000110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011110011001100110011001100110111011101110111101110111011101110111011011101110111011101110111011101110011001100110011001100110010111011101110111011101110111011101110111011101110111010101010101010101010101010101110111011101110111011110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100110001000100001000100010010001000100100100010011001100110011001,
	2400'b100110011001100110101010101010101010101010101010101010101001100110000111011001100111100010011010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111011111111111011101111111011101110111111101111111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011011101110111001011101110101010101010011001100110011000100010001000011101110111011101110111011101110111011101110111011101100110011001100111011101110111011101111000101010101001011101100110011101110111011101110111011101111000100010000111011101110111100010001000100001110111011101110111011101100111011101110111011101110111011101110111011101110111100010001001100110011000100010011011110011001100110011001100101110111010101010101010101010111011101110101010101010010011000100010010001000100111110011001100110011001100110011011100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111100110011001100110011011101110111011101110111101110111011101110111011101101110111011101110111011100110011001100110011001100101110111011101010101010101010101010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001000100001000100010010001000110100100010011001100110011001,
	2400'b100110101001100110101010101010101010101010101010101010011000100001110111100010001001100110011001101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111001100110011001100110010111011101110111011101110111011101110111010101010101001100110011001100010001000100001110111011101100110011001100110011001110111100001110110011001100111011101110111011101110111011101110111100001110111011101110111100010001000011101110111011001100110011001100110011001100110011101110110011101110111011101110111011101111000100001110111011110001001101010111011101110111011101110101001100110011001100110101010101010101010101010100100000100010001001000100110101110111011101110111011101110111011101010101010101010101010101010101011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110111011101110111101110111011101110111011011101110111011101110111011101110111011101110111001100110011001100110011001100110010111011101110111011101110111011101010101011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011010101010100110001000100001000100010010001000110100100010011001100110011001,
	2400'b101010101010101010101010101010101010101010101010101010101001100110011001100110011010100110011010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110101011101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110011001100110011001100101110111011101110111011101110111011101110111011101110111010101010101001011101100110011001100101011001100110011001100110011001100110011001100110011001100110011001110111011101110111011001100111011101110110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111100010011010100110101010100110000111011110001000100010001000100110011001100110010011000100100010001000100101101010101010101010101001100110011001100110001000100010001000100010001001100110011010101010111011101110111011101110111011110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011100110011001011101110111011101110111011101110111011101110111011101110101010101010101010101010101011101110111011101110111011101110111011101110111011110011001100101110111011101110111011101110101011101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001101010100110001000100001000100100010001000100100100010011001100110011001,
	2400'b101010101010101010101010101010101010101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111110111011101111111111101110111111111110111111111111111111111110111111101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100101111001100110011001100101110111011101110111010011101100101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101100110010101100110011001100110011101110111011110000111011101111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010000011001000100010001000100100100110011001100110011001100110001000100010001000100001110111011101110111011110001000100110101010101110111011101110111011101111001100110011001100110011001100110011001100110011011101110111011101110010111011101110111010101010101010101110111011101110111010101010101011101110111100110011011101110111011101110111011101110111011101110011001100110010111011101110111011101110111011101010101010101010101010101010011010101010011010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010100110001000100001000100100010001000110101100010011001100110011001,
	2400'b101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011101101111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011011100110011001101110011001100101110111011101110100111011001010101011001100110011001100110011001100101010101010101010101010101010101010101011001100110011001100110011001010101010101010101010101010101010101010101010101010110011001100111011101110111011101110111100110101010101110111011101010101001100001110111011101110111011101110111011101111000100010001000100010001000100010001000100010000100000100100010001000100100100110011001100110011001100010001000100010001000011101110111011101110111100010001000100010001001100110111100110011001100110011001100110011001100110011001100110011001101110111011101110111001011101110101010101010101010101010101010101010111011101010101001100110011001100110011010101010111011101111001100110111011101110111011101110111001100101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101001100110011010101010101011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010100101001000100001000100100010001000110101100010011001100110011001,
	2400'b101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101010101010100110011010101010111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111011101110111111101110111111101110111111101110111011101110111011101110111011101110111011101110111111101110111011101110111011101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110010111011101110111011101010010111011101110111011101110111011101110111011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011101110111011110001001101010101001100110111100101110101000011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010000101001000100001000100100011100010011001100110011001100010001000100010001000100010000111011101110111011101111000100010001000100110101010101111001100110011001100110011001100110011001100110011001101110111011101110011001011101110111010101010101010101010101010101110111011101110111010101010011001100110011001100110011001101010101010101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101111001100110011001011101110111011101110111011101110111011101110111011110011001100110011001100110011001011101110111011101110111011101110111011101110111010101010100101001000100001000100100010001101000101100010011001100110011001,
	2400'b101010111011101110101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101010101010100110011001101010111011101110111011101110111011101110111011101110111011101110101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101110111011101110111111111111111111111110111111101110111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101010101010100101110110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001010110011001100110011110011001100001110110011110011011101110000111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010000101001000100001000100100011100010011001100110011001100110011001100110001000100001110111011101110111011101110111011110001000100010001000100110011001101010111100110011001100110011001100110011001100110111011100110011001011101110111010101010101010101010101011101110111011101110111011101010101010101010011001100110011001100110011001100110101010101010111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011100110010111011101110111011101110111011101110111011101110111100110011001100110010111100101110111011101110111011101110111011101110111011101110111010101010100101001000010001000100100010001101000101100010101001101010011001,
	2400'b101010111011101110101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001101110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111111101110111111111110111111111111111111111111111111111110111111101110111011111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110111011101110111001100110011011101110111011101110111011100110011001100110011001100110011001100101110111010100110000111011101110110011001100101010101010101010101010101010101010101010101010101010101010101010101010101011001100110010101010101010101010110011101110110011001100110011010001010100101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010000101001000100010001000100011100010011001100110011001100110001000100010001000100010001000100001110111011101110111100010001000100010001000100010001000100010011001100110011001101010101010101010101010101010111010101010101010101010101010101010101010101010101010101110111011101110111011101110101010101010101010101010011001100110011001100110011001100110101010101010101011101110111011101110111011101110111011101110111011110011001101110111001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010100101001000010001000100100011001100110100100010101001101010101001,
	2400'b101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001101110111011101110111011100110011001100110011001100110011001100110011001100101110111010100101110111011001100110011001100101010101010101010101010101010101010101010101010101011001100101010101010101010101100111011001010110011001100110011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000110001000100001000100100010011110001000100010001000100010001000100010001000100010001000100010001000100010001000100110101001100110001000100010001000100010001000100010001000100010001000100010011001100110011001100110011010101010101010101010101010101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101011101110111011110011011100110011001100101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010100101001000010001001000100010001100110100100010101010101010101010,
	2400'b101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100101110101001100110001000100001110111011101100110011001100110011001100110010101010101010101010101010101010101011001110111010101010110011001100110011001110111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110101001000010001000100100010011010001000100010001000100010000111011110001000100010001000100010001000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001101010101011101110111011101110111011101110111011101110111011101110101011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101010101010101110111010101010100101000100010001000100100010001000110100100110101010101010101010,
	2400'b101010101010101010101010101010101001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011100110011001100110111001100110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100110011001100110011001100101110111010101010101010101010011001100110011000100010001000011101110110011001010110011001110111011101110110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110101001000010001000100100010010110000111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001101010111011101110111011110011001100110010111011101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111010101110101010101010101010101010101010101010101010101010100101000100010001000100010001001000100100100110111010101010101010,
	2400'b101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110101001100010001000100010001000100110011001101010101001100001110110010101010110011001100110011001100110011001010110011001010101010101010101011001100110011001100110011001100110011001100111011101111000011110000111011110000110001000100001000100100001010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001101010101010101110111011101010011001100110011001100110011010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100000100010001000100010001001000110100100110111010101010101010,
	2400'b101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011101111111111111111111111111111111111111111111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100110011001100110011001100110011001100110011001100101110111011101110111011101010011001100110011010101010011001100110001000100010000111011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001110111011101110111011101110101001000010001000100100010010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110101001100110011001100110001000100010001001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010100000100010001000100010001001000110100101010101010101010101010,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110010101000100010001000100010001000011001100110011001101000100010101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001001100010001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001000100010001000100010001000011001100110011001100110100010001010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100001110111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101110111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110011001100110011001100101010101000100010001000100001100110011001100110100010001010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100010001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100001110111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010111011101110101010101110111011101110101010101010101010101010101010101010101010101010101010101110111011101111001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100010001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110010101010101010101010101010101010100010001000100010000110011001100110011010001010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100001110111011101111000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010011001100110011001100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010100110011010101010111010101010101011101110111011101110111011101110111011101110111010101010101010101110111011101010101010101010101011101110111011110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110010101010101010101010101010001000100010001000100010000110011001100110011010001010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010001000100010011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011101110111011101110111011110001000100010001000100010001000100010011001100110011001100010011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100110011001100110011000100010001000100010001000100010011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110100010101101000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110011001100110010101010100010001000100010001000100001100110011001000110011010001010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010001001100110001000100110011000100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000111011101110111011101110111011101110111011101110111011110001000100010001000100010011001100110011000100010011001100110011001100110011001100110011001100110011001100010001000100010001001100110011001100110011001100110011000100010001000100010001000100010011001100110011001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011110000111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110100011010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011101110111011101100101010001000100010001000100001100110011001100110011010001010111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110001001100110001000100010001001100110011001100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100110001000100110011001100110011000100010001000100010001000100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001101010111100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001100111011101100110011001010100010000110011001100110011001100110011001101010111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011000100110001000100110001000100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011000100010001000100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101001100110101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011110001000100001111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001000110011001100110100011110001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011001100110011001100101010000110011001100110011001100110011001101010111011101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010000111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010011001100110001001100110011001101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101111001011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100010011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010000111100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001100110011001101101000100010001000100001111000100010001000100010001000100010001000100010001000011101110110011001010101010101100101010101000011001100110011001100110011001101000110010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111100110010111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001100100010001000110101100010001000011101100111011110001000100010001000100010001000100010001000100001110111011101100101010101010101010101010100001100110011001100110011001101000100010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011000100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001001100010011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001001100110011001100110011010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001100110010001100110011010101111000100001100110011101111000100010001000100010001000100010001000100010001000011101100110010101010100010101010100010000110011001000110011001101000100010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011000100010011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011001100110011001101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110011001100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111100001111000100010001000100001110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111,
	2400'b010000110011001100110011001100110011001100110011001101000110100001100101011001100111100010001000100010001000100010001000100010000111011101110110010101010100010001000100010000110011001100110011001101000100010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011000100110011001100110011001100110001001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011000100010011001100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100001111000100010001000100010001000011101110111100001110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101000100010001000011001100110011001100110011001100110011010101100100010101010110100010001000100010001000100010000111100001110111011101100110011001010101010001000100001100110011001100110011001100110100010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001111000100001111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101010101000100001100110011001100110011001000110011001101000100010001010101011001110111100010001000100010000111011101110110011001100110011001010101010001000100001100110011001100110011001100110100010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011110001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100001111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101010101000100001100110011001100110011001100110011001100110011010001000101010101100111100010000111011101110111011101110110011001010101010101100101010001000100001100110011001100110010001100110100010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100010001001100110011001100110011010101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010000111011110001000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101100101010001000101010000110100001100110011001100110010001000110011001100110100010001010110011101110111011110000111011101100110010101010101010101010101010101000100001100110011001100110010001000110100010001010110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011010100110101010101010011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110010111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100001111000100010001000100001111000100010000111100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010100010001000100010001010101010001000011001100110011001000100011001100110011010001010101011001111000011101110111011101100110010101010100010101010101010101010100001100110011001100110011001000110011010001010101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001101010101010101010101010101010101010101010101010101010011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001011110010111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001110111100001111000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101000100010001000101011001100110010101010100010000110011001000110011001100110011001101000101010101010111011101110111011101100110010101010101010001000100010001010101010000110011001100100011001100100011001101010101011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011110010111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101111000100001111000100001111000100010000111100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101010101000101010101010100010001000100010001000011001000100010001000100011001101000100010001010110011001110111011101100110011001010100010001000100010001000100010000110011001100110011001100100011001101000101011001010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011000100110011000100010001000100010001000100110011001100110011001100110011001100110011001100110001001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100001110111011110000111011101110111100010000111011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101000100010001000100001100110011001100100010001100110011001100100010001000100010001100110011001101000101010101110111011101110110011001100101010001000100001100110011010001000011001000110011001100110010001101000101010101000110011110001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110001000100010011001100110011000100010011001100110011001100110011001100110011001100110011000100110001001100110011000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111100110011001011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011110000111011101110111011101110111011101110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101011001100101010001000011001100100010001000100011001100100010001000100010001000110011001101000100010101010110011001110111011001010101010101000011001100110011001100110100001000100011001100110010001001000100010101010110011110001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010011000100110011001100110011001100110001001100010001001100110011001100110011001100010011000100110011001100110011001100110001001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011110011001011101110111100101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101110111011101110111011110000111100001110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101100110010101010101010000110011001000100010001000100010001100110010001000100011001100110011010001000101011001100110011001100101010101010100001100110011001100110011001100110011001100110010001000110100010101010110011001111000100010001000100010001000100010001000100010001000100001111000011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010011001100010001001100110011001100110011001100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111100110011001100101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110110011001010100010001000101010101010100001100100010001000100010001000110011001100100010001100110011010001000100010101010101010101100110010101000100010000110010001000100011001100110011001100110010001000110100010001010101011001111000011110001000100010001000100010001000100010001000011101100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100101010101010100010001000100010101010100001100110010001000100010001000110011001100110010001000110011001100110011010001000100010101010101010101010100001101000011001000100010001100110011001100100010001000110100010001010101011001100111011110001000100010001000100010001000100010001000011001000101010101010110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110010101010100010001000100010001000100010000110011001000100010001000100011001100110011001000110011001100110011001100110100010001000100010001000100010000110011001100100010001000110010001100100010001000110100010001000101010101100111100010000111100010001000100010001000100001110110010101000100010001000100011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110010101010101010101010101010001000100010001000011001100100010000100100010001100110011001100100011001100110011001100110011001100110100010001000100001100110011001100110010001000100010001000100010001000110100010001000100010101010111011101111000100010001000100010000111011101100101001100110011001101000110011001110111011110001000100010001000100010001000100010001000100010001000011101100111011101111000011101110111100010001000100010001000100010001000100010001000100010001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110010101010101010101010101010101010101010101000011001100100010000100010010001000110011001100100011001100110011001100110011001100110011010000110100001100110011001000110011001000100010001000100010001000110100010001000100010101010111011101110111011110000111011101110110011001010011001100100011010001000100010001000101010101100111011110001000100010001000100010001000100010000110010101100111011101100110011001100111011110001000100010001000100010001000100010001000100110001000100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011001100110010101010100010001000100010000110011001100100010001000100010001000100010001100100010001000110011001100110011001100110011010000110011001100110011001100100011001100100010001000100010001000110100010001000100010001010110011110000111011101110111011101100101010000110011001000100011001101000100010001000100010101010101010101100111011110001000100010001000011101010110011101110111011001100110011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110111011101110111011101110111011101110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110011001100110011001100101010101000011001100110011001000100010001000100001000100100010001000100010001000100011001100110010001100110011001100110011001100110011001000100010001000110010001000100010001000110011010000110100010001010101011101110111011001100110011001000100001100110011001100110011010001000100010001000100010001000101010101010110011001100111011101110110010001100111011101010101011001100110010101010101010001000100010001000100010001010110011101111000100010001000100010001001100010001000100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011110111011101110111011101110111011101101110111011100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101100110011001010101010001000011001100100010001100100010001000010001000100010011001000100010001000100011001100110011001000110011001100110011001100110011001000100010001000100011001000100010001000110011010000110011010101000101010101100111010101100100010000110011001100100011001101000100010001000100010001000100010001000101010101010101010101010101010101000011010101100100001100110100001100110011001100110011001100110100010001000100010001000100010001010101011110001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111100010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110110011001100101010101000100001100100010001000100010001000100001000100010010001100100010001000100010001100100011001100110011001100100100010000110011001000100010001000100010001000100010001000100011010000110100001100110101010101100101010101000011001100110011001100110011010001000011010001000100010001000100010101010101010101010101010101000100001100100011001100110010001000110011001100110100010001000100010001000011010001000100010001000100010001000101010101010111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110110111001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100010001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101111000011101110111011001100110010101010100010000110010001000100010001000100010001000010010001000110011001000100010001000110010001000100011001100110011001100110011001000100010001000100010001000100001001000100011001100110100001000110100010101010100001100110011001100100010001100110011001101000100010001000101010101010100010101010101010101010100010000110010001000100010001000100011001101000100010000110011010001010100010001000100010001000100010001000100010001000100010101010110011110001000100010001000100010001000100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111011110011001100110011001100110011001100110011001100110011001100110011001100110111101110111011101110111011101110111011101110111011101110111011101110111011011101110011001100110011001100110011001100110011001100110010111011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b100010001000011101110111011001100101010101000100010001000011001100100010000100010001001000100010001000110011001100100010001000110011001000100010001000110011001000100011001000100010001000100010001000100001001000100011001100110011001100110011010001000011001100110010001000100011001100110011001101000100010001010101010101010101010101010100010000110011001000100010001000100010001000110011010001000100010101010100001101000100010101000100010101010110011001010100010001000100010001000101011001111000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111011101111001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001100110011001011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101110111011101110110011001100110011001010101010001000100001100110010001000010001000100010001001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110010001100110011001100110100010001000100010001010100010001000100010101000100001100100010001000100010001000100010001100110011001101000100010001000101010001000100010001010100010001100111011101110110010101010101010001000100010001010110100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001011101111001100110011001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110111001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101111000011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001001000110011101110110011001010101010101010101010101000100010000110011001000010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010000100100010001000010010001000100010001000100010001100100010001000100010001100110010001000100011001100110011001100110100010001000100010001010101010001000100010000110010001000100010001000100010001000100010001000110011010001000100010101000100010001000100010001000101010001010110011110001000011101100101010101000100010001000100011110001000100010001000100010001000100010001000100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110111101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011001110111,
	2400'b000100100011010001100111011101100101010101010101010101000100010000110011001100100010000100010001000100010010001000100010001000100011001000100010001000100010001000100001000100010010001000100010001000100010000100100010001000100010001000100010001000110010001000100010001000110011001100110100010001000100010001010101010001000011001000100010001000100010001000100010001100110011001100110011001101000100010001010101010101010100010001000101010101010101011001111000100001110110010101010101010001000100010101111000100010001000100010001000100010001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011001110110011101100110011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110,
	2400'b000100010001001001000101011001100101010101010101010101010100010001000011001100100010001000010001000100010001001000100010001000100011001100100010001000100010001000100010000100010001001000010010000100010001001000100010001000100010001000100010001000100010001000100011001100110011001100110011001101000101010101000100010000110010001000100010001000100010001000100010001100110011001100110011001100110011010001000101010101010101010001000100010101010101010101111000100010001000011101100101010101000100010001011000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101100111011001110110011001100110011101110110011101110111011101100111011101110111011101110111011101110110011101110111011101110111011101100110,
	2400'b000100010001001000100011010001010110011001010100010101010100010000110011010000110010001000010001000100010001000100100010001000100010001100110010001000100001001000100010001000010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001100110011001100110100010001000100010001000100001100100010001000100010001000100011001100110010001100110100001100110011001100110100010001000101010101100101010101000100010101100101010101010111100010001000100001110101010101000100010001000110100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110110011001110110011001100110011101100110011101100110011101100110011101110111011101110111011101110111011101110111011101110110011101110111,
	2400'b000100010001000100010001001000100100010101010101010101000100010000110011001100110010001000010001000100010001000100010010001000100010001000110011001000010001000100100010000100010001000100010001000100010010000100100010001000100010001000100010001000100010001000100010001000110011001100110100001101000100010001000010001000100010001000100011001100110011001100110011001100110011010001000100010001000100010001000100010101100110010101010100010101100111011001010110100010001000100010000111011001010100010001000100011010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001110111011101110110011001100110011001100110011001100110011001100110011001110110011001110111011101110111011101110111011101110111011101110111011001110111,
	2400'b001000100001000100010001000100010010001101000101010001000100010001000011001100110010001000100001000100010001000100010001001000100010001000110011001000010001000100010001001000010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110010001000100010001000100010001100110011001100110011001100110011001101000100010101000100010001000100010101010110010101010101010101010111011101010101011110001000100010001000100001100100010101000100010001111000100010001000100010001000100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101111001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011101110110011001110110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011001110111011101110111011101110111,
	2400'b001000100010000100010001000100010001001000110010001101000100010001000011001100110011001000100010000100010001000100010001000100100010001000110010001100100001000100010001000100100001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001000100010001000100010001000110011001100110011001100110011001100110011001101000100010001010101010101010101010101010101010101100110010101010110100001110110010110001000100010001000100010000110011001100101010001010111100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110110011101110110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000010001000100010001001000100001001000100010001100110011001100110011001100110011001000100001000100010001000100010010001000100010001100110001000100010001000100010010000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001000100011001100110011001100110011010000110011010001000100010001010110011001010110010101100101011001100111011001010101011110000111011001111000100010001000100010001000011110000110010101000101100010001000100010001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110011001100110011101110110011001100110011001100110011001100110011001100110011001100111011001110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100010001000100010001000100010001000100010001000100100010001100110011010001000100001100100001000100010001000100010010001000100010001100100010000100010001000100010001001000010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001000100010001100110011001100110011001100110011010001000011001101000100010101010101011101100110011001100110010101110111011001100101011001110111011101111000100010001000100010001000100010001000011001010100011010001000100110011000100010011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100111011101100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001001100110011010000110011001000100010001000010001000100010001000100010010001000100010001000010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001100100010001000010010001000100010001000100010001000100011001100110011010001000011001101000011001100110101010001010101011010000111011101110110011001111000011101110110011001100111011110000111100010001000100010001000100010001000100001110110010110001000100010001000100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011101110110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100100100010000110011001100100001000100010001000100010001000100010001000100010010001000010001000100010001000100010010000100010001001000010010001000100001000100010001001000100010001000010001001000100010001000100010001000100010001000100010001000100010001000100011001100110011010001000100001100110100010001000100010101010101011001111000100001110111011101101000100001110111011001100111100010001000011110001000100010001000100010001000100010001000011001111000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011101110110011001100110011001100110011001100101011001100110011001100111011101100111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010010001000100001000100010001001000100001000100010010001100110011001000100010000100010001000100010001000100010001000100010001000100100001000100010001000100010001000100010001001000100001001000010010001000100010001000100010001000010001001000100010001000100001001000100010001000100010001000100010001000110011001100110011010001000100010001000100010001000100010101010110010101100111100010000111100001111000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111100010001000100010011001100110011001100110011001100110011001100110011000100010011000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011001100110011101110110011001100110011001010101010101000101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010001000100010010000100010001000100010001000100010001000100100011001000100001000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100010001000100010001000100100010001000100001000100010001000100010010001000100010001000010010001000100010001000100010001000100010001000110010001000110011010001000100010001000100010001010101010101100110011001100110011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000111011101110111100010011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011001100110011101110110011001100110010101010100010001010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100100010000100010001000100010001000100010001001000010001000100010010001000100010001000100010001000100010001000110011001100110011010001000100010001010100010001000101010101010110011001100110011001111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001110111011101110111011101110111011110001001100110011000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010000111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011001110111011001100110011001100110011001100101010000110100010101010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100100001000100010001000100010001000100100010000100010001000100010001000100100010001000100010001000100010001000100010001000100011001100110011001101000100010001010101010101100101011001110110011101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011110001001100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101110110011001100110011001100011001101000101010101010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000010001000100010001001000100010001000100010001000100010001100110010001000100011001100110011010001000100010001010101010101010110011001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010001000100010001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111011101110111011101110111011101110111011110001000100010001000011101110111011110000111011110001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001110111011101100101010100110011001101000100010101010101010101010110011001100111011101110111011101110111011101110111011101110111011101110111011001110111,
	2400'b001000110010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001101000100010101010101011001010101011101110111100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001101111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001110111011101110111011101110111011101110111100010001000100001110111011001110111011101110111011101111000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110110011001100110011001000100010000110011010001000100010101010101010101010110011001110111011101110111011101110111011101110111011101110111011101110111011001110110,
	2400'b001100110010001100100010001000010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001100110010001000100010001000100010001000100010001100100010001100110011001100110011010000110100010101010101011001100101011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110111101111111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101001100110011001100110011001100110011001100110011000100010011001100110011001100110011001100110011000011101110111011101110111011101110111011101111000100010001000011101110111011101110111011101110111011101110111100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011101100101001100110010001100110100010001000100010001010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110110,
	2400'b010000110100001100110010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100011001000110010001000110011001100110100010001000100010001100101011001110111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110111011110111011101110111011101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011000100010011001100110000111011110001000100110011001100110001001100110001000011101110111011101110111011101110111011101111000100010000111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011101010011001000100010001000110101010001000100010001010101010101100110011001100110011101110111011001110111011101110111011101110111011101110111011101100110,
	2400'b010001010101010001000100010000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100100001000100010001000100100001000100100010001000100001001000100010001000100010001000100011001100110011001000110011001100110011010101010101010001000110011001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011011101111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110011001100110000111011110001000100001110111011101111000100110011001100010001000100010000111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111100010001000100010001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110010100110011001100100010001000110101010001000100010001010101010101100110011001100110011001100110011001100111011101110111011101110111011101110111011101100110,
	2400'b010001100101010101010101010100110010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000010010001000010001001000100010001000100010001000100011001100110011001100110011001100110011010001010110010101010101011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011000100010001001100110001000100010001000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100111011101111111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001011101110111011101110111011101110111011101111000100010011001100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110010000110010001100110010001101000100010001000100010001010101010101010110011001100111011101100110011001110110011001110111011101110111011101110111011101100110,
	2400'b011001100101011001100110010000100011001100100010001000100001001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000010001000100100001000100010001000100010001000100100001001000100010001000010001000100100010001000100010001000110010001101000011010001000011001100110011001101010110011001100101011001110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010011001100010011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011011110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011000011101110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100110011101100101001100110010001100110010001101010100010001000100010001010101010101010110011001110111011101100110011001100110011001110111011101110111011101100110011001100110,
	2400'b011001100110011001100101001100110100001100100011001100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100010001000100010001000100010010001000100010001000100010000100010001001000100010001000100010001000110011001000110100001101000100010101000011001101000110011101100110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010011000100010011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001101111011101110111111111110111011101110111111101110111011011100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100101110111011101110111011101110111011101110111011101111000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011001100100001100110010001100110010001101010101001101000100010001000100010101100110011001110110011101100110011001100110011001110111011101110111011101100110011001100110,
	2400'b010101010110011001100101001101000100001001000100001100110011001000010010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100001001000010001001000100010001000100010001100100011001100110011010000110011011001010011010001000110011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011011110111011111111111111111111111011101101110111001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100001110111011101110111011101110111011101110111011101111000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110110011001100101001100110011001100100010001101000101010001000100010001000101011001100110011001100110011001100110011101100110011001110111011101100110011001100110011001100110,
	2400'b010101010101010101010011001101000011001101010100001101000011001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100001001000100010001000100010001000100010001100110011010001000011001101000100010101100100010001000101011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111100110011001100110011001100110011001100110011001100110111011101111011011101110111001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011000011101110111011101110111011101110111011101110111011101111000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001110111011101110111011101110111011101110111011101100111011101110111011101110110010101010100001100100011001100100010001101000101001101000100010001000101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001010101010101000100010001000011010001000100010001000011001000110011000100010001000100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010000100100010001000100010001000100010001000100010001000110011001100110011001101000100010001010101010001010101010101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101001100110011000011101110111011101110111011101110111011101110111011101110111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101011001110110011101110111011001110111011101110111011001110110011001100110011001100110010101010100001100110010001100110010001101000101010001000100010001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001010101010101010101010001000100010001000100010000110011001100110010000100010001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100010001000100100010001000100010001000100010001000100010001000100011001100110100010001000101010001000101010101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101010101010101100110011001110111011101100111011101110111011001100110011001100110011001100101010101000100001100110010001100110010001101000101010001000100010001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b010101010101011001010101010101000100010001000100001101000100001100110011001000010010001000010010000100010010000100010010001000010001000100010001000100010001000100010001001000100001000100010001000100010001000100010001000100010001001000100001000100010001000100010001000100010010000100010010001000100010001000100010001000100010001000100011001100110100010001000101010101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100110011001100110011001010101010101010110011001110111011001100110011001100110011001100110011001100110011001100101010101000100001100110010001100110011001101000100010001000100010001000101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b001000100011001100110100010101010100010001010100010001000011001101000011001100110010001000010001000100100010001000010001000100010001000100010001000100010001000100010001001000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100001001000100010001000100010001000100010001000110011001101000100010001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110101001100110101001100110011001100110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110011001100110011001010100010001010101011001100110011001100110011001100110011001100110011001100110011001100101010001000100001100110010001100100011001101000100010001000100010001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100010010001100100010001000110011001100110100010001000100010000110010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100100011001100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100100001001000100010001000100010001000100010001000110011001100110011001101000100010101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100010000111100010011001100110011010100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110010101010101010001000101010101100110011001100110011001100110011001100110011001100110010101010101010001000011001100110011001000100010001101000011010001000100010001010101010101010101010101100110011001100110011001100110011001100101010101010101011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100100011010001000100010100110011001100100010001000110011001000100001000100100001000100010001000100010001001000100001000100100100010000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010010001000100010001000100010001000100010001000110011001100110011001100110011001100110100010001010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110000111011101110111100010011001100110011001100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101011001100110011001010101010101000100010101010110011001100110011001100110011001100110011001100110010101010101010001000011001100110010001100110010001101000011001101000100010101000101010101000101011001100110011001100110011001010101010101010101010101010110011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100010001001000110011001100110011001100110011001100110100001100100010001000100010001000100010000100010010001000110011000100010010010000110001001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010010000100010010001000100010001000100010001000100010001100110010001100110011001100110011001100110011001100110011010001010110011110001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100001110111011101110111100110011001100110011001100110011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101011001100101010101000011010001010101011001100110011001100110011001100110011001100101010101010101010000110011001100100010001100110011010000110011010001000100010001000101010001000101010101100110011001100110010101010101010101010101011001100110011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001001000100011001100110011010000110011001100100010001000100010001000100010001000010001001101000100001000010001001100100001001101000010001100100001001000010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001101000011001100110011010000110100010001010110100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001110111011101110111100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001011101110111011101111000100110011001100110011001100110011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101010101010101010101010100001101000110011001100110011001100110011001100110011001010101010101010100010001000011001100110010001000110011010001000011010001000100010001000100010001010101010101100110011001100101010101010101010101100101011001100110011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011001100110011001100100010001100110010001100110011001100110001001001000100001100010001001000010001001100110011001000010010001000010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001100110010001100110011001100110011001100110011001100110011001100110100010001000100010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100001110111011101110111011110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000011101110111011101111000100010001000100110011001100110011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010001000101010001000101010001000101010101100110011001100110011001100101010101010101010101000100001100110011001100110011001000100011010001000011001101000100010001000100010101010101011001100110011001010101010101000101010101010110011001100110011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100011001100100010001100110011001101000100010000110011000100110100001100100001000100010001001100110010001000100010000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011010000110011001100110011001100110100010001000100010001000101011001100111100010001000100010001000100010001000100010001000100010011000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110011000100010001000100010001000100010001000011101110111011101110111011101111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010111011101110111011101110111011101111000100110011001100110011000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101000100010101000100010000110100010101010110011001100110011001100110010101000100010001000100001100110011001100110011001000110011010000110011001101000100010001000101010101010101011001100110010101010101010001010101010101010101010101100110011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001100110011010000110101010101000100001000100100001100010001000100010001001000100001001000100001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011010001000100010001000011010000110011010001000100001100110100011001100101010101000101010101100111100010001000100010001000100010001000100010001000100010001000100010001000100110001000100110011001100110011001100110011001100010011001100010011001100110011001100110011001100110011000100010001000100010000111100010000111011101110111011101111000100001110111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000111011101110111011101110111011101110111100110011001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101010011010001010100010001000011010001000110011001100110011001100101010101000100010001000100001100110011001100110011001100110011010000110011001101000100010001000101010101010110011001100101010101000100010001010101010101010101010101100110011001100110011001100110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001100110011001100110011010101010100001100010010010000100001000100010001001000010001001000010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001000100010001000100010101010100010001000100010001000100001101000100010001100111011101100101010001000101011001111000100010001000100010001000100010001000100010001000100010001000100110001000100010001001100010001000100010001000100010001000100010001000100010011001100110011001100110011000100010001000011101110111011101110111011101110111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110010111011101110111011101110111011101110111100110011001100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101010100001101000100001101000011001101000101011001100110011001100101010101000100010001000011001100110011001100100010001000100011010000110011001101000100010001010100010101010110011001010101010001000100010001000100010001010101010101100110011001100110011001100110,
	2400'b001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100011001001000011001101000101010000100001001100110001000100010001001000010010001000010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000110010001000110011001100110100010001000100010001010101010101010101010001000100010001000100010001000100010001000101011001110111011001010100010101010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000100010001000011101110111011101110111011101110111011101110111011110000111011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110000111011101110111011101110111011101111000100110011000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100101010101010101010000110011010001000011001001000100011001100110011001100101010101010100001101000011001100110011001100100010001000100011010000110011010001000100010001000100010101010101010101010100010001000100010001000100010001010101010101100110011001100110011001100110,
	2400'b001000100001000100010001000100010001001000100001001000010001000100010001000100010001000100010001000100100010001000110010001100100010001000110101010000110100010000110001001000110001000100010001000100010011001000010001000100010001000100010001001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001000100010101010101010101010101010101000100010001010100010001000100010001000100010101100111011101110110010101010101011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100001110111011101111000011101110111011101110111011101110111011101111000011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100001110111011101110111011101110111100010001000100110011000011110001000011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010100010101000011001100110011001000110100010101100110011001100101010101010100010000110011001100110010001000100010001000100011010000110011010001000100010001000101010101010101010101000100001101000011001100110011010001010101010101100110011001100110011001100101,
	2400'b001000100010000100100010001000010010001000100010001000100010001000100010001000100010001000010010001000100010001000100011001101000011000100010010001101000011010000110001000100100001000100010001000100100011000100010001000100010001000100100011010001000010001000100010001100100010001000100010001000100010001000100010001000100010001000110010001100110011001100110100010001010101010101010101010101000100010101010101010101000100010001000100010001000101011001111000011101100101010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001111000011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110000111011110001000011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010001000100010000110011001000100011010001010110011001100101010101010100010001000011001100110011001000100010001000110100010000110011010001000100010001000100010101010101010001000100001100110011001100110011010001000101010101100110011001100110011001010101,
	2400'b001000100010001000100010001000100010001100110011001100100011001100100010001000110010001000010011010000110011001101000011001100110100010000100001000100110011001000100001000100100001000100010001000100100010000100010001000100010010001000110010001000100010001000110011001100110010001000100010001100100010001000100010001000100010001100110010001100110011001100110011001100110100010001010101010101010101010101010101010101010100010001000101010101010101010101100111100001110111011001010101010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100001110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010101000011010000110011001100100010010001010110011001100101010101000100010001000011001100110011001000100010001000110011010000110011001100110100010001000100010001010100010001000011001100110011001100110100010001010101011001100110011001100110011001010101,
	2400'b001000100010001100110010001000100011010001010101001100100011001100110010001100110010001000010011010101000100010001010100011001010100010001000100001000010001001000010001000100010001000100010001000100100001000100010001000100010010001000100010001000110011010001000011001101000011001000110011001100110011001100100010001100110010001000100011001100110010001100110010001100110011001100110011010000110100010001010101010101010101010101010101011001100111011001010111100001111000011101110101010001010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100001110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101010100001100110011001100100010001101000101010101100101010001000100010000110011001100110011001000100010001000110011010000110011001100110100010001000100010001000100010000110011001100110011001101000100010101010110011001100110011001100110010101010101,
	2400'b001000110011010000110010001000110100011001100100001001000100001100110011001100100011001000100100010101000110010101100110011001110110010101010100010000100001000100010001000100010001000100010001000100010001000100010001000100010001001101000100010001000100010001000011010001000011001100110011001100110011001100100011001100110011001100110011001100110011001100100010001000110011001100110011001100110011001100110100010001010101010101100101011001100111011001000110011110001000011101110111011001010100010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101111000100010011001100110011001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011000011101110111011101110111011101110111011101110111011101110111011110001000100010001001100110011001100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101100110011001100110011001100111011101100111011101110110011001100110011001010101010101000100010001000011001100110010001000110101010101010101010001000011001100110011001100110011001000100010001000110011001100110011001101000100010001000100010000110100001100110011001100110011010001000101010101100110011001100110011001100101010101100101,
	2400'b001001000110010100100011001100110101010101010011010001000011001101000011001100110010000100100101010101010110011001100110011001100110011001100110011001000010000100010001000100010001000100010001000100010001000100010001000100010100010101100101010000110100010001000100010000110010001000110010001101000100001100110011010001000100001101000100010001000011010000110011001100110011001100110011001100100011001100110011001100110100010101010101010101010101010001000100011001110111011101110111100001110110010101010110100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110011001100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100010000111011101110111011101110111011101110111011101110111011101110111100010001000100110011001100110011001100110011001100010001000100010000111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010100010000110011010001000100010000110011010001000100010101010110011001100110011101110110011001100110010101010101010001000100010001000011001000100010001000100100010101010101010101000100001100110011001100110011001000100010001000100011001100110011001100110011001101000100001101000011001100110011001100110100010101010110011001100110011001100110011001010101011001100101,
	2400'b010001100111010000110101010001010110011101010100011001010100010000110011010000110001000100110101010001100110011001100110011001100110011001100110010101000010000100010001000100010001000100010001000100010001000100010001000100010011010101100110010101000100010101000100001100110010001100100010001101000100001100110011010001010100001101000100010001000100010101000011010001000011001100110011001100100011001100110011001100110011010001000100010101010101010101010101010101110111011110001000100010000111011101100101011010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011110001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111100010001001100110001000100110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110001000011101110111011101110111011101110111011101110111011101110111011110001000100010001001100110011001100110011001100110011001100110011000100010000111011110001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010001000011001100110011001100100010001000100010001000100010001000100011001101000100010101100110011001100110011001100101010101000100010001000100010001000100001100100010001000100011010101010100010001010100001100110011001000100011001000100010001000100011001100110011001100110011010001000011010000110011001100110011010001000100010101010101011001100110011001100110010101010101011001100101,
	2400'b011101110110010001100101010001100111011101000110011001010101010000110011001100100001000100110100010001010101010101010101010101000100010000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110010001000100010001000100010001000110011001101000100001100110011010001010101001101000100010101010100010101010100010001010100010001000100001100110011001100110011001100110011001100110011010001010101010101010101010101100111011110001000100010001000100001110111010101111000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001111000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000100001110111011101110111011101110111011101110111011101110111011101110111100010001000100010011001100110011001100110011001100110011001100110011000100010001000011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101000100001100110011010001000100001100110011001000110010001000100010001000100011001100110011001101000101011001100110011001100101010101010100010001000100010001000100001100100010001000100011010001010100001100110100001100110011001000100010001000100010001000110100001100110011001100110011001100110011010000110011001100110011010001000100010001010101011001100110011001100101010101010110011001010101,
	2400'b011101110100010101010101010101100111011001100111011001010100001100110010001000010001000100100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100011001100110011001101010101001101010101010101010100010101010100010101010100001101000100010000110011001100110011001100110011001100110011010001000100010101010101011001100110011110001000100010001000100001110111011101110111100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011110001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111100010001000100010000111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001000100001110111011101110111011101110111011101110111011101110111011101111000100010001001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010001000011001101000100010001000011001100110011001100110011001000100010001000100010001000100010001000110011001101000101011001100101010101010100010001000100010000110100001100110010001000100010010001000100001100110011001100110010001000100010001000100010001000110100001100110011001100110011001100110011010001000011001100110011001101000100010101010101011001100110011001100101010101100110011001100110,
	2400'b011001010110010101010101010101110111011001110101010100110011001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000110100001101010101011001100101011001100100010101010100010001000100001101000100010001000011001100110011001100110011001100110100010001010101011001100111011110001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101100111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100010001000011101110111011101110111011101110111011101110111011101110111011101111000100010001001100110001000100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100001110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010101000100010001000100010001000011001100110011001100100010001000100010001000100010001000100010001000100010001000110011010001010110010101010101010001000100001101000100010000110011001000100010001101000100001100110011001000110011001000100010001000100010001000110100001100100011001100110011001100110011001100110011001100110011001101000100010101010110011001100110010101010101011001100110011001100110,
	2400'b010101100110010101110110011101100110010101010100001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000110100010101100101011001100101011001010101010101000100010001000100010001000100010001000011001100110011001100110100010001000101011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001100110011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100010001000011101110111011101110111011101110111011101110111011101110111011101111000100010001001100110001000100010011001100110011001100110011001100110011001100110001000100010001000100001111000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101100110010001010101010101000100010001000011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001100110100010101100101010101000100010000110100001100110011001100100010001001000011001100100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011010001000100010101010101010101100101010001010110011001100110011001100110,
	2400'b011001100110011101110110010101010100001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010001000100100010001000100010001000100010001000100010001000100010001000110100010101010101011001100101011001010101010101000100010001000100010001000100010000110011001100110011001101000100010101100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101100101010101110111011001100110011110001001100110011001100110000111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011110001000100010011001100110011000100010011001100110011001100110011001100110011001100110011000100010011000100010001000100010001000100010001000100001110111100001110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101011001100101011001100101010101000101010001000011010000110011001100110011001100110011001100100010001000100010001000100010001000100010001000100010001101000101010101000100010000110011001100110011001100100010001000110011001000100010001000100010001000100010001000100010001000100010001100110011001000110011001100110011001100110011001100110011010001000101010101010110011001100101010001100110011001100110011001100110,
	2400'b011001010110011101010101001100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110100010101100101011001100101011001010100010001000101010101010101010101000100001100110011001101000100010001010111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011001010101010101100110011001100110011110001001100110011001011101100110011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011000100110011000100001110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100110011000100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100001110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010110011001100110010101010101010101000100010001010100001100110100010001000100010000110011001100100010001000100010001000100010001000100010001000100011010101010100010000110011001101000011001100100010001000110011001000100010001000100010001000100010001000100010001000100010001000110011001000110011001100110011001100110011001100110100010001000101010101010101011001010100010101100110011001100110011001100110,
	2400'b011001010100001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100001000100010010000100010001001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100011001101000101011001100110011001100101010101000101010101010101010101010100010100110011001100110011001100110110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101110110010101010101010101100101011001100110011110001000100110000111011001100110011001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110001000100010001000011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110001000100110011000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101100110010101010110010101010101010101010100010001010100010001010101010001000100001100110010001000100010001000100010001000100010001000100010001101000100010001000011001100110011001100100010001000110011001000100010001000100010001000100010001000100010001000100011001000100010001000110010001000110011001100110011001100110100010001010101010101010101010101000101011001100110011001100110011001100101,
	2400'b010000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001000100010000100010010000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011010001010101011001100101010101010101011001010110011001100101010101010100001100110011001100110100011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011001100110011001100110010101010110011101110111011101110111011101100101010101010101010101010101011001100110011110001001100001100110011001100110011010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110101010101010011000100010001000100010000111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110001001100110011000100010001000100010001000100010001000100010000111011101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110010101100110011001100110011001100110010101010101010101010101010101000100010000110011001100100010001000100010000100010001000100010001001000100011010001000011001100110011001100100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000110011001000110011001100110100010001010101010101010101010001000101011001100110011001100110010101010110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100011010000110010001100100010001000010010001000100010001000110011001100110011001100100010001000100010001000100010001000100010001000110011001101000100010001010101011001100101011001100110011001100101011001100101010000110011001100110011010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011001110111011001100110011001100110011001010110011001110111011101110111011101110101010101010101010101010101011001100111100010001000011001100110011001100110011001111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011010100110001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100110011001100110011001100110011001100110011000100010011001100110001000100110001000100010001000100010001000100010001000100001110111011001100110011001100110011001100110011101110111011001100110011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110110011101110110011001100110011001010100010001000100001100110011001100100010001000100010000100010001000100010001000100010001001000110011001100110011001100100010000100100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001100110011001101000100010001000101010101010100010001010110011001100110011001000100010101100110,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010010001000100010010001000100010001000011001100110010001000100010001000110100001100110011001100110010001000100010001000100010001000100010001000100011001101000100010001000100010101010110011001100110011001100110011001110110010100110100010000110011001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011001110111011001100110011001100110011001010101011001110111011101110111011101110110010101010101010101010101011001100111100010000110011001100110011001100110011001111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010101010101001100110011000100010001001100110011001100110001000100010001000100001111000100001110111011101110111011101110111011101111000011101111000100010001000100010001000100010001000100010001000100010001001100110011001100110011000100010011001100110011000100010011000100010001000100010001000100010001000011101110111011001100110011001100110011001100110011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101100110011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011001100110011001100110011001000011001100110011001100110011001000100010001000100010001000010010000100010001000100010001000100010011010000110011001100100010000100100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001000101010101000100010101010110011001100100001000110101010101010101,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000010001000100010010001001000100010001010101001100110100001100110011001100110100010001000100001100110011001100100010001000100010001000100010001000100011001100110011010001000100010001010101010101100110011001100110011001110110011001000100010001000011001101000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100110011001100110011001100110011001010101010101100111011101110111011101110101010101010101010101010101011001100111011101100110011001100110011001100111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011000100010001000100010011001100010001000100010001000100010001000100001111000100001110111011101111000011110001000100010001000100010001000100010001000100010001000100010011000100010001000100010001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110011001100110011001010101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101000100010001000100010000110011001000100010001000110011001000100010000100010010000100010001000100010001001100110011001100110010000100100010001000100010001000010010001000100010001000100010001000110011001000100010001000100010001000100010001000110011001100110100010001010101010001000101010101100110010000100011010101100110011001010100,
	2400'b000100010001000100010001000100010001000100010001000100010001001000010001000100010010000100010010001000110010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100001000100010010001000100011010001010110011000110101010101000100010001000100010001000100010000110011001100100011001000100011001100110011001000110011001100110011001101000100010001010101010101010101011001100111011001110110011001100100010001010011001100110100011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001010101010101100110011001100110011101100101010101010110011101110111011101110110010101000101010001010101011001110111011001010101011001100110011001111000011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110001000100010001000100010001000100010011001100010001000100010001000100010000111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110011001100110010101000100010001000100011001110111011101110111011101110111011101110111011101110111011101110111011001010110011001000101010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100101010001000100010001000100001100110011001000110011001100100010001000100010001000100001000100010001000100010001000100100010001100100010000100010001001000100010001000100010001000100010001000100010001000110011001000100010001000100010001000100010001000110011001101000100010001000100010001000101011001100011001000110101010101100110011001000011,
	2400'b000100010001000100010001000100010001001000010001000100010010001000100001001000100010000100010010001000100011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010000100010010001000100010001101000110011001100100010001010100010001000100010001000100010001000011001100100011001100100010001000110011001100110011001100110011010001000100010001000100010101010101011001100111011001110111011001100110010001010100001100110011010001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011001100101010101010101010101010101011001100110010101010101011001110111011101110101010001000100010001010101011001100110010101010110011001100110011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100010001000100010001000100010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011001100101010001000011001100110011010001010110011001100110011001110111011101110111011101110111011101100110010101010101010101010101010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101010101010101000100010000110011001101000011001100100010001000100010001000100001000100010001000100010001000100010001001000100010000100010001001000100001000100100010001000100001001000100001001000110011001000100010001000100010001000100010001100110011001101000100010001000011001101000110010100100011010001010110010101100101010000110011,
	2400'b000100010001000100010001000100010001000100010001001000010010001000100010001000100010001000100010001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010000100010010001100110100010101100110001100110100010101010101010101010101010101000011001100110100010000110010001000100010001100110011001100110011001101000100010001000100010001000101010101100110011101110111011101100110010001000100001100110011001101000110100010001000100010000111100001110111100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110011001100101010101010101010101010101010101010110010101010101010101100111011101110101010101000100010001000101010101010101010101010101010101100111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000100010001000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100101010001000011001100110011001100110101011001010110011101100110011001110111011101110111011001010101010001010100010001010101010101010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011001010101010001010101010001000100001100110011010001000011001100110011001000100010001000010001000100010001000100010001000100010001000100010010000100010001000100010001000100010010000100010001000100010001001000100010001000100010001000100010001000100010001100110011001100110100010000110011010001010100001000110101010101100101010101010100010000110010,
	2400'b000100010001000100010001000100010001000100100010001000100010001000100010001000100011001000100010001100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010000100010010001100110011001101000100010101000100010001000100010001010101010101010100010000110100010101000010001000100010001100110011001100110011001100110100010001000100010001000100010101010110011001110111011101100111010101000100001100110100001100110100011101110111011101110111011101110111100010001000100010001000100010001000100001110111100010001000100001110111011101110111011101100110011001100110011001010101010101010101010101010101010001010101010101010110011101100110010101010100010001000101010101010101010001000101010101010111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100010000111011101110111100010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110010101010100010001000100001100110011001100110100011001010101011001100101011001100110011101110110010101000100010001000100010001000100010001000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101010101010101010101010101000100010001000100001101000011001100110010001000100010001000010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000110010001000100010001000100010001000100010001100100011001100110011001000110101010100110010010001010101011001010100010001010011001100110010,
	2400'b000100010001000100010001001000100001001000100010001000100010001000100011001000110011001000100010001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100100010001000100010001000010010001000100100010000110011001100110100010001000100010001000101010101010100010001000100010101000011001100110011001100110011001100110011001100110100010001000100010001000100010001000101011001110111011001110111011001010100001101000100010000110011010101110111011101110111011101110111100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101100110011001100110011001100101010101010101010101010100010001000100010101010110011001100110010101000100010001000101010101010101010101000101010101110111011101111000100010011001100110011001100110011001100110011001100110011001100110011000100010001000100010001001100110011001100110011001100110011001100110001000100001111000100110011001100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010011000011101110111011101110111011101111000100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001100110011000100010001001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110010101010101010001000100001100110011001100110011010001010100010101010101010101100110011101100101010001000011001100110100010001000100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101010101000100010001000100010001000100001100110011001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000110010001000100010001000100010001000100011001100110011001100110010001101010101001100100101010101010101010101000011001100110011001000100010,
	2400'b000100100010001000010010001000100010001000110010001000100011001100110011001100110011001000100011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010010001000011001100110010001000100010000100010011001101000011001100100011010001000100010001000101010101010101010101010100011001010100001100110011001100110011001100100011001100110011010001000100010001010101010101010101010101110111011101110111011001010101010001010100010001000011001101010110011101110111011101110111011101110111011110001000100010001000100010000111011101110111011101110111011101110111011101100110011001100110011001100110010101010101010101010100010001000100010001010101010101100101010101000100010001000100010001010101010001000101010101100110010101010110011101110111100010001001100110011001100110011001100110011001100110011000100010001000100010001000100110011001100110011001100110001000011101110111011101110111100010011001100110011001100110011001100110011001100110001000100010001000100010011001100110011001100110011010101010101010101010101010101010101010101010101010101010101001100110000111011101110111011101110111011101110111011101111000100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001111000100010001000100010001000100010001000011101110111011101110110011001100101010101000100001100110011001100110010001101000011001101000100010101010110011001010100001100110011001100110011001100110100010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101010101010101010101000101010001000101010101000100010000110010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100011001100110011001100110100010101010100010001010101010101010011001000100010001000100010001000100010,
	2400'b000100010001000100010010001000100010001000110011001100100011001100110100001100110011001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010001010100001100110011001000100010001000010010001100110100010000110011001100110011010001000101010101010101010101100101010101100101001101000011001100110011001100100011001100110011010001000100010101010101010101010101010101100111011101110111011101100101010101010101010001000011001100110101011001110111011101110111011101110111011101110111100010001000100010001000011101110111011101110111011101110111011101110110011101110111011101100110011001100101010101010100010001000100010001000100010101010100010001000100010001000011010001000100010101010101010101010101010101010110011001010101011001111000100010001001100110011001100110011001100110011000100010001000100010001001100110011001100110011001100010000111011101110111011101110111011110001001100110011001100110011001100110011001100001110111011101110111011110001000100110011001100110011001100110101010101010101010101010101010101010101010101010011000011101110111011101110111011101110111011101110111011101110111100010001001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010000111011101110111011101110110011001010101010001000100010000110011001100110010001000110010001100110100010001010101011001010100001100110011001100110011001101000100010101010110011101110111011101110111011101110111011101100111011001100110011101110111011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101100101010101010101010101010100010001000101010000110010001100110010001000100010000100100001000100010001000100010001000100010001000100010001000100010001000100100001000100010001000100010001001000100010001000100010001000100010001000100010001100110011001001000101010101000100010101010101010000110010001000100010001000100010001000100011,
	2400'b001000100010001000100010001000110010001000110011001100100011001101000100010000110011001100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001010101001100110100001100100010000100010010001000110100010001000100001100110010001000110100010101010101010101100101010101100101001101000011010000110011001100110011001100110011001101000100010101010101010101010101011001100110011101110111011101110110011001010110011001010100010001000100011001110111011101110111011101110111011101110111011110001000100010001000100010000111011101110111011101110111011101110111011101110111011001110111011001100110011001010101010001000100010001000100010001000011001100110100010001000100010001000100010001000100010101010101010101010101010101010101011001100110100010001000100110011001100110011001100110011000100010001000100010001001100110011001100110001000100001110111011101110111011101110111011101111000100110011001100110011001100110011000011101110111011101110111011101110111100010001001100110011001101010011001100110011010101010101001101010011001100110000111011101110111011101110111011101110111011101110111011101110111011101111000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110110011001100110010101000011001100110011001100100010001000100010001000110011001101000101011001010100001100110011001100110011010001000100010101010110011101110111011101110111011101110111011001100110010101100111011101110111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001010101010101010100010101010101010000110011001100110011001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100001000100010010001000100010001000100010001000100010001101000101010101010101010101010100001000100010001000100010001000100010001000100010,
	2400'b001000100010001100100010001100110011001000110011001100100100010001000101010100110011001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001010110011001000100010100110010001000010001000100100100010101010101010000110011001100110011010001010101011001100110011001100110010001000100010000110011001100110011001000100011001101000100010001010101010101010101011001100110011001100111011101110110011101100110011001100100010001100100010001100111011101110111011101110111011101110111011101110111011110001000100010001000011101110111011101110111011110001000011101110111011001110111011001100110011001100110011001000100010001000100010001010100001100110100010001000100010001000100010001000101010101010110010101010101010101010101011001100110011010001000100010001000100010011001100110011000100010001000100010001000100110011000100001110111011101110111011101110111011101110111011101111000100110011001100110011001100110000111011101110111011101110111011101110111011110001001100110011001100110011001101010101001100110011001100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101111000100110011010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000100001110111011101110111011101100110010101010100001100100010001100100010001000100010001000100011001101000101010101000100010000110011001100110011001101000100010101100110011101110111011101110111011101100110010101010101010101100110011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100101010101010101010101010101010001000100001100110011001000100011001100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100110010000100100010001000100010001000100010001000100011010001000101010001010101010000100010001000100010001000100010001000100010001000100010,
	2400'b001000100011001100110010001101000011001000110011001100110100010101000101010000110011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001010110011001010100010001000010001000100010001000100011010001010101010000110011010000110011001000110101011001100110011001110110010001010100010001000011001100110011001000100010001100110100010001010101010101010110011001100110011001100111011101110111011101110110011101100110010001100110010101010110011101110111011101110111011101110111011101110111011101110111100010001000011101110111011101110111011110000111011101100110011001100110011001100110011001100110011001100100010000110100010001000101001100110100001101000100010001000100010001000100010001010110010101010101010101010101010101010101011001111000100010001000100010001001100110001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010011001100110011001100001110111011101110111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001101010011001100110101001101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000011110001000100010001000100010001000100001110111011101110111011101100110010101010101010000100010001000100010001000100010001000100010001100110100010001000011001100100010001100110011001101000100010101100110011101100111011101110111011001010101010001010101010101100110011001110111011101110111011101110111011101100110011101100110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011001110111011101110111011001100101010101010100010101010101010001000011001100110011001100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000110100010001000100010000110010001000010010000100100010001000100010001000100010001000100010,
	2400'b001000110011001100110011010001000100001100110011010000110100010101010100001101000011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001010101011001100110010001000011001000100010001000100010001101010101010101010011010001000011001000110100010101010110011001110110010001100101010001000100001100110011001000110011001100110011010001000101010101010110011001100110011001110111011101110111011101110111011101110111010101010110011001010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101100110011001100110011001100110010101010101010101100101010000110100010001000100010000110011001101000100010001000100010001000100010001000101010101010101010101010110011001010101011001111000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111100010001001100110011000100001110111011101110111011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111011110001001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000011101100110011001010101010101010110011001111000100010001000100010001000100010001000100001110111011101110111011001100110011001100101010100110010001000100010001000100010001000100010001000100011010001000100001100100010001100110011001101000100010101010110011001100110011101100110010101000100010001000101010101010110011101110111011101110111011101110110011001110110011001110110011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011001100110011001010101010001010101010101000011010001010100001100100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000110011001100110010000100010001000100010001000100010010001000100010001000100010001000100010,
	2400'b001100110011010001000100001101010101010000110100010001000101010101000011010001000011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001000101010101100111011001000011001000100010001000100010001000110101010101010100001101000101001100110011001101010110011001110110010101010101010001000100010001000011001100100011001100110011001101000100010001010110011001100110011001110111011101110111011101110111011101110111011001100110011001100101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100101010101010101010101010101010101000100010001000100010000110011001100110100010001000100010001000100010001000101010101010101010101010110011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011101110111011101110111011101110111011110001000100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100110101010100110011001100110011001100110101010100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010000111011001010101010101000100010001000100010001010110011110001000100010001000100010001000100010000111011101110110011001100110011001100101010001000100001100100010001000100010001000100010001000100011001101000011001100110011001100110011001101000100010001010101010101100110011001100101010101000100010001000100010101100111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010101010101010001000101010101000100001100110010000100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001100110010001000010001000100010001000100100001000100010001001000100010001000100010001000100010,
	2400'b001100110011010001000100010001010101010000110101010101000101010001000101010000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100100011010001000101010101100111011001100011001000100010000100010010001000100100010101000101010000110100010101000011001101000101011001100110011001100100010101010100010001000011001100110011001100110011001100110100010101010101010101100110011001110111011101110111011101110111011101110111011101110111011101100110011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010101010101000100010001000100010101010100010000110100010001000100010001000100010001000100010001000100010001000101010101010101010101010110011001100110011001100111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011010100110011001100110011001100110011010100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100001110101010101000100010001000100010000110011001101000100010101100111100010001000100010001000100010001000011101110110011101100110011001100101010101010100001100100010001100100010001000100010001000100011001100110011001000110011001100110011001101000100010001010101010101100110011001010100010001000100010001000100010101100110011101110111011101110110011001100110011001010101010101000100010001000100010101010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011001100110011001110110011001100110011001100101010001010101010101000011010000110010001000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100010010001000100001000100010001000100010001000100010001001000100001000100010001001000100010001000100010,
	2400'b001100110100010001000100010001010110010000110110011001000100010001010100010000110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000010001000100010001000100100011010001010101010101100111011001100101001100100010001000100010001000100010010001010101010101000011010001000011001100110100010001010110011001100110010101010100010001000011001100110011001000100011001100110011010001010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101100101010101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100110011001100110011001100101010101010101010001000100010001000100010001000100001100110011001100110011001100110011001101000100010001000100010101000101011001010110011001100110011001100110011101100111100010001000100010000111100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000011101100110011001010101010101000100010001000100010001000101011001111000100010001000100010000111011101110111011001100110011001010101010001000100001100110011001000110010001000100010001100110011001100110010001000100011001100110011001100110011010001010101010101010101010101000100010001000100010001000100010101010110011101110111011001100110011001010101010001000100010001000100010001000101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100101010101010101010001000100010000110011001100100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010000100100010000100010001000100010001000100010001000100010001000100100010001000010010001000100010001000100010,
	2400'b010001000100010001000101010101100110010101000110011001000101010101010100010000110011000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100010001001000010001000100010001000100010011010001010101010101100110011001100101010000100010001000100010001000100010001001000110010101010011010001010100001100110011010001000101011001110111010101010101010101010100010001000011001000110011001100110011010001010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110110010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001010101010101010101010101010101010001010100010001000100001101000100001100110011010000110011001101000100010001000101010001000100011001100110011001110111011101110111011101111000100010001000100001110111011101111000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100110011001100110011001100110011001100110011001100110011001100110011000011110001000100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100101010101000100010001000100010000110011010001010110011110001000100010000111011101110111011001100110011001010101010101000100001100110011001000100011001000100010001000100010001100110010001000100011001000110011001100110011010001010101010101010101010101000100010000110100010001000100010101100111011101110110011001100110010101000100010000110100010000110011010001000100010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011101100110010101000100010001000011010000110011001100100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001100100010,
	2400'b010001000100010101010101010101100110010101000110010101000101010001000100001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100010001000100010100010001010101011001100110011001010101010000110010001000100010001000100010001000110100010101100101001101010101010000110011001101000100010001100111011001100101010101010101010000110011001100110011001100110011010001000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011001110110010101100101010101010101010101010101010101000100010001000100001100110100001100110011001100110011010001000100010001000101010101010101010101100111011101110111100010001000100010001000100010001000100010000111011101110111100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100110011001100110011001100110011001100110001000100010000111011101110111100010000111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001010101010001000100010001000100010001000100010001100111100001111000100001110111011001100101010101010101010101000011001100110011001000100010001100100010001000100010001000100010001000100010001000100010001100110011010001000100010101010100010001010100010001000100010001000101011001100111011001100110011001010100001100110011001100110011010001000100010001010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101100110011001100110011001100110011001100110011001100110011001100110010101010100010001000100001100110011001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001001000010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000110011,
	2400'b010001010101010101010101011001100111010101010110011001000101010001000011001100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000010001000100010010000100010001000100100100010101010110011001100110011001010101010000110010001000100010000100100010001000100011010001100110010001000101010101000011001100110011010001010111011101100110010101010101010001000100001100110011001100110011001100110100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010110011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100110011001100110011001100110011001010101010101010100010001000011001100110011001101000100001100110100010001000011010001000100010101010101010101010111100010001000100010001000100010001000100010001000100010001000011101110111100010011000100110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010011001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100110010101010101010001000100010001000100010001000101011110001000100001110111011101100101011001010101010001000100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010001000011010001000100010001000100010001000101011001100110011001100101010000110011001100110011010001000100010001010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100110011001100110011001100110011001100110011001100110011001100101010101010100010101000100010000110011001100100010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100001000100010001000100010001000100010010000100010001000100010001001000100010001000110011001000110011,
	2400'b010001010101011001100110011001110111010101010110010101000101010000110010001000010001000100010001000100010001000100010001000100010001000100010001000100100010000100010010001000100010000100010001000100010001000100110101010101010110011001100110011001010101010001000011001000010010001000100010000100100010001101000110010101000101010101010100010001000100010001010110011101110111011001100101010101000100001100110011001100110011001100110100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101100110011101110111011101110111011101110111011101100111011001100110011001100110011001100101010101010101010101010100010001000100001100110100001100110100001100110011001100110011001101000011010001000100010001010110011110001000100010001000100010001000100010001000100010001000100010001000100010011000100010000111011101110111011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110011000011110001001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001001100110011001100110000111011101110111011101110111011101110111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001010101010101000100010001000100010001000101010101100111100001110111011101100101010101010101010101000100010000110010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010000110011001101000101010101000100010101100110010101000011001100110011001101000100010101010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010100001100110011001000100011001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100100011001100110011001000100001000100100010000100010001000100010010001000100010001000100010001000100010001000100011001100110011,
	2400'b010001100101011001100110011001110111010001010110010101000100001100110010000100010001000100010001000100010001000100010001000100010001000100010001001000100010000100010010001000010010000100010001000100010010001000110101010101100110011001100110011001010101010001000011001000100010001000010010001000100010001000110101011001000101010101010101010001000100010001000101011001110111011001100110011001010101001100110011001100110011001100110011010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110110011001110111011101110111011101100111011101110110010101100110011001100110011001100101010101010100010101000100010001000011001100110011001100110011001100110011001100110011001100110011010001000100010001000101011001111000100010001000100010001000100010001000100010001000100010001000100010001001100010000111011101110111011001100111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100110000111011101111000100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101111000100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100101010101000101010101000100001101000100010001000101011001110111011101110110011001010101010001000011001100100010001000100010001000100010001000100010001000100010001000100011001000100010001000110011001101000011001100110011001100110011010001010101010101000101011001010100001100110011001100110011001101000100010001010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111011001110110011001100110011001100110011001100110011001100110010101100110011001100101010101010100001100110011010001000011001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110100010001000100001100100001000100010001000100010001000100010001001000100010001000100010001000100010001100110011001100110011,
	2400'b010101100101011001100110011101110110010001100110010101000011001100100001000100010001000100010001000100010001001000010001000100010010000100010001000100100001000100010001001000100001001000010010000100010010001101000101011001100110011001100110011001010101010101000100001000100010000100010010001000010001001000100011010101100100010101000101010101000100010001000100010101100111011101100110011001010101010000110011001100110011001100110011010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110110011101100110011101110111011101110111011101100110011101100110011001100110011001100110011001100110010101010101010001000100010001000011010001000011001100110011001100110011001100110100001100110011010001000100010001000101010101100111011101110111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110011001100111011101100110011001100111011101110110011101110111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100001110111011101110111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101111000100010011001011101110111011101110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100110010101010101010101010100010001000100010001000100010001100111011101110110011001010101010000110011001000100010001000100010001000100001001000100010001000100010001000100010001000110010001000110011001100110011001100110011001100110100010001000101010101010101010000110011001000100010001000110011001101000100010101010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101110110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010001000100001100110011001100110010001000010001000100010001000100010001000100010001000100010001000100010001000100010001001001000101010001000011001000010001000100010001000100010001000100100010001000100010001100110011001100110011001100110011001100110011,
	2400'b010101100110011101100110011101110110010001100110010000110011001000010001000100010001000100010001000100010001001000010001001000100010001000010001000100100001000100010001000100100010001000010001000100010010010101100110011001100110011001100110011001000101010001010101001000110010001000100001001000100001001000100010001101100110010101100101011001010100010001000100010001010111011101110110011101100110010001000011001100110011001100110100010001010111011101110111011101110111011101110111011101110111011101110111011101100110011101100110011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110110011001100110011001100110011001100110010101010100010001000100010001000100010000110011001100110011001100110011001101000100010001000100010001000100010001000100010101100111011101110111011101110111011101111000100010001000100010001000100010001000011101110111011001100110011101100110011001100111011001110110011101100110011001110111011001110111011101110111011101110111011110001001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110011001100110010101010101010001000100010000110100010001000101011101110110011001010101010101000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001101000100010001010101010101000011001100110010001000100010001000100011001100110011010001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101100110011001100110011001100110011001100110011001100110011001100110010101010101010001000100010001000100001101000100001100110010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001101010101010000110010000100010001000100010001000100010001000100100010001000100011001100110011010001000011001100110011001100110011,
	2400'b010101100110011101110110011101110101010001100110001100110011000100010001000100010001000100010001000100010001001000100001001000100010001000010001000100100001000100010001000100010010001000100010001000100100011001100110011001100110011001100110010101010101010001010101001100110010001000100010001000100010001000100010001000110101011001100101011001010101010001000100010001010110011101110111011101110110010101000011010000110011001100110100010001100110011101110111011101110111011101110111011101110111011101110111011101100110011101110110011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110110011001100110011001100110011001100110010101010100010001000101010101010100010001000100001100110011001100110011001100110100010001000100010001000100010001000100010001010110011001100111011101110111011101110111011101111000100010001000100010000111011101110111011101110110011001100110011001100111011001100110011001100110011001100110011101110111011101110111011101110111011110001001100110011001100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110011001110110011001010101010101000100010000110011010001000101010101100110011001010110011001010011001000100010001000100010001000100010001000100010001000100010001100100010001000100010001100100011001100110010001100110011010000110100010101010101010000110011001100100010001000100010001000110011001101000100010101010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100101010101010101010001010101010101000100010001000100010001000011001100110010001000100010000100010001000100010001000100010001000100010001000100010001000100010011010001000100001100100001000100010001000100010001000100010001000100100010001000110100010001000100010001000100010001000100010001000011,
	2400'b010101100111011101110111011101110101010101100100001100100001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100001000100010010001000010001000100100010001000100101011001100110011001100110011001100110010101010101010101100101010000110010001100110010001000100010001000100010001000100011010101100110010101100101010101000100010001000101011001110111011101110111011001010100010101000011001100110011010001010111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101110111011101110111011101110111011101110111011001100111011101110111011101110111011001100110011001100110011001100110011001100101010101000100010001010101010101010101010001000100001100110011001100110011001100110011010001010100010001000100010001000100010001010110011001100110011001110111011101110111011101110111100010001000100001110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011110001001100110001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001100110011001010101010101010101010001000100010000110011010001010110011001100110010101010100001100100010001000100010001000100010001000100010001000100010001100110011001000100010001000100011001100110011001100110100001100110101010101000100001100110010001000100010001000100011001100110100010001010101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001010101010101000101010101010101010101010101010101000011001100110011001100110010001000010001000100010010000100010001000100010001000100010001000100010001000100100100010101000100001000010001000100010001000100010001000100010001001000100011001100110100010101000100010001000100010001000100010001000100,
	2400'b011001100111011101110111011101110100011001100100001100010001000100010001000100010001000100010010001000010010001000100010001000100010001000100010001000100001000100010001001000100010001000010001001001000110011001100110011001100110011001100110011001010101011001100101010000110011010001000010001000100001001000100010001000100010001101010110010101100110010101010100010001000101011001110111011101110111011001100101010101000100001100110011010001010110011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100101010001000100010101000101010101010100010001000100001100110011001100110011001100110011010001010101010001010100010001010100010001010101011001100111011101110111011101110111011101110111011101111000100001110111011101110111011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111100010001001100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001100110010101010110010101010101010101000100010001000011001101000101011001100110010101010101010000110010001000100010001000010010001000100010001000100010001000110010001100100010001000100010001000110011001100110011010001000100010001000011001000100010001000100010001000100011001100110100010001000101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110110011001100110011001100110011001100110010101010101010101010101010101010101010101010100010001000100001100110011001100100010001000100010001000100010001000010001000100010001000100010001000100010001001001000101010101000010000100010001000100010001000100010001000100010010001000110011010001000100010101010011010001000100010001000100010001000100,
	2400'b011001100111011101110111011101100100011001010011001000010001000100010001000100010001000100100010001000010010001000100010001100110010001000110010001000010001000100010001000100010001001000100001001001010110011001100110011001100110011001100110011001100110011001100101001100110011010001000100001000100001000100100010001000100010001000110110011001100110011001010100010001010101010101100111011101110111011001100110011001010100010001000011010001010110011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011001100110011101100100010101010101010101010101010101000100010001000011001100110011001100110011001100110011010001000101010101010101010101010101010001010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011110001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001010110011001100110010101010110010101010101010101010100001100110011010001010101010101010101010101000011001000100010001000100010001000100010001000100010001000100010001100100010001000100010001100110010001100110011010001000100010000110010001000100010001000100010001000110011001101000100010001000101010101010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011001100110011001100110011001100110011001100101010101010101010101010101010001000100010001000100010001000011001100110100001100100011001100110010001100100010001000100010001000100010000100010001000100010001000100110100001100110010000100100001000100010001000100010001000100100010001101000011001100110011001100110011010000110011001100110100010001000100,
	2400'b011001100111011101110111011101000101010100110010000100010001000100010001000100010001000100010001000100100010001000100010001101000011001100110010001000010001000100100001000100010001000100010010001101010110011001100110011001100110011001100110011001100110011001100101001100110100010101000100001000100010000100100001001000100010001000100011011001110110011101100101010001000101010101100111011101110111011101100110011001010100010001000011001101000110011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011001100101011001100110010101010101010001000100010001000011001101000011001100110011001100110011001100110100010101010110010101010101010101010101011001100110011001100111011101110111011101110111011101110111011101110111011001100111011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100111011101100101011001100110011001100110011001010100010000110011001101000101010101000100010001000011001000100010001000100010001000100010001000100010001000100010001100100010001000100010001100110010001100110011010001000100001100100010001000100010001000100010001100110100010001000100010001010101010101010101010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100110011001100110011001100101010101010101010101010101010101000100010001000100010001000011010000110011001100110011001101000011001100110010001100110011001100110010000100010001001000100001000100110011001100110001001000010001000100010001000100010001001000100011001100110010001000100010001000100011001100110011001100110011001100110011,
	2400'b011001110111011101110111011001000101010000100001000100010001000100010001000100010001000100010001000100100010001000100010001101000100001100110010001000010001000100010001001000100010001000010010010101100110011001100110011001100110011001100110011001100110011001100101010001000101010101010100001000100010001000100001001000100010001000100010010001110110011001100101010101010101010101010110011101110111011101100111011101100101010001000100001101000101011001110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110110011101110111011101110111011101110111011101110110011101100110011001100110011001100101010101000100010000110011001100110011001100110011001100110011001100110011001100110100010001010110011001010110011001010101011001100110011001100111011101110111011101110111011101110111011101110111011001110111011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001110111011101100111011101100110011101110110011001010101010101000011001100110100010101000011001101000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000011001000100010001000100010001000100010001100110011001100110100010001000101010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110010101010101010101010100010001000100010001000011001100110011001100110011001100110011001100110011001100110010001000110011001000100010000100010001001000100001000100100010001100100001001000010001000100010001000100100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011,
	2400'b011001110111011101110111010101000100001100010001000100010001000100010001000100010001001000010001001000100010001000100010001100110100001100110010000100010001000100010001000100010001000100100100011001100110011001100110011001100111011001100110011001100110011001100101010101010101010101010101001100100010001000100001001000100010001000100010001101010111011001100101010101010101010101010110011101110111011101110111011101100110010101010100001100110101011001110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101110111011101110111011101110111011101110110011001100110011001100100010001000100010000110011010000110011001100110011001100110011001100110011001100110100010001000101011001100110011001100101011001100110011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111100010001001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011001110111011101100110011001100110010101010101010001000100001100110011001101000011001100110010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100011001100100011001100110010001000100010001000100010001000100010001000110011001100110100010001010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011001100110011001100110011001100110011001010101010101010100010001000100010001000100001100110011001100110011001100110011001100100010001000100010000100010001000100010001000100010001000100100001000100100011001000010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000110010001100110010001100110011,
	2400'b011101110111011101110110010001000011001000010001000100010001000100010001000100010010001000010010001000100010001000100010001100110100001100100011001000010001000100010010001000100001000100100101011001100110011001100110011001100111011001100110011001100110011001100110010101100110011001100101001100110010001000100010000100010010001000100010001000110110011101100110010101010101010101010110011101110111011101110111011101110110010101010101010000110100011001110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011001100110011001100110011001010100010001000100010001000100010000110011001100110011001100110011001100110011001100110100010001000100010101100110011101100101011001100110011001110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110110011001100110010101010100010001000100001100110010001000110100001100100010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001100110100001100100010001000100010001000100010001000100011001100110011001101000100010001000101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101100110011001100110011001100110011001010100010001000100010001000100010001000100010001000100001101000011001100110011001100110010001000100001000100010001000100010001000100010001000100010001000100100010001000010001000100010001000100010010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011,
	2400'b011101110111011001010100001100110010001000010001000100010001000100010001000100010010001000100010001000100010001000100010001101000100001100100011001000010001000100010001000100100001000100110110011001100110011001110111011101110111011101110110011101100110011001100110011001100110011001100101010000110010001000100010001000100010001000100010001000110100011001100110011001010101011001100110011101110111011101110111011101110111011001010110010101000100010101100111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101100110011001100110010101010100010001000100010001000101010000110011001100110011001100110011001100110011010000110011010001000100010001010110011001100110011001100110011101100110011101110111011001110111011101110111011101100110011001110110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001001100110011001100110011001100110011000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101100101010101010100010001000100001100110010001100110011001100110010001000100010000100100010001000010010001000100001000100100010001000100010001000100010001000100010001100110011001000100010001000100010001000100010001100110011001100110011001100110100010001000100010101010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110111011001100111011001100110011001100110011001100110011001010101010001000101010101000100010001000100010001000100010001000011001100110011001100100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001100110011001100110011010000110011010000110100,
	2400'b011001100101010001000100001000100010000100010001000100010001000100010001000100010010001000100010001000100010001000100010001101000100010000110011001000010001001000010001000100100010001001000110011001100110011101110111011101110111011101110111011001100110011101110110011001100110011001100101010001000011001000100010001000100010001000100010001000100011010001100110011001100110010101100110011001110111011101110111011101110111011101100110010101000100010001100110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011001100110011001100101010001010100010001000100010101100101001100110011001100110011001100110011001100110011001101000100010000110100010001010110011001100110011001100110011001100110011101110111011101110111011101110111011101100111011101100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011110000111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100001110111011101100110010101010100010001000100010000110011001100110011001100110010001000100010000100100010000100100010000100010001000100100001001000100010001000100010001000100010001100110010001000100010001000100010001000100010001000100010001000110011010001000100010001000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110010101000101010101000100001100110011001100110011001100100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100011001100110011001100110011010001000100,
	2400'b010001000100010001000011001000100010000100010001000100010001000100100001000100100010001000100010001000110011001000100010001101000100010000110011001000010001000100100001000100010001001001000110011001100111011101110111011101110111011101110111011001100111011101110110011001100110011001100101010101000011001000100010001000100001001000100010001000100010001101000101010101100110011001100101011001110111011101110111011101110111011101100111011001010100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011001100111011001100100010001000100010001000101010101010100001100110011001100110011001100110011001100110011001101000100010001000100010001000101011001100110011001100110011001100110011001100111011001100111011101100111011101110111011001100110011101100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111011110001000100010000111011110001000011101111000100001110111011101100101010101010101010001000100010000110011001100110011001100100010001000100010000100010001000100010010001000010010001000100010001000100010001000100010001000100010001100100010001000100010001000100010001000100010001000100011001100110011010001000100010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011001100110011001100110011001100110011001100110011001100110011001100101010101000011001100110010001000100010001000100010001000100001001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001100110011001101000100010001000100010001000100,
	2400'b010001000100010001000010000100100010000100010001000100010001000100100001000100100010001000100010001000110011001000110010001001000100010001000011001000010001000100100010001000010001001001010111011001100111011101110111011101110111011101110111011101110111011101100110011001100110011001100101010101010011001000100010001000100010001000100010001000100010001000110100010101100110010101100101011001110110011101110111011101110111011101110111011101010100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011001100110011001110111011101110111011101110111011101110111011001100110011001010100010001000100010101010101011001010100001100110100001100110011001100110011001100110011001101000100010001000100010001000100011001100110011001100110011001100110011101100111011101100110011101110111011001100110011001110110011001100110011001100110011001100110011001100110011001100110011101100110011101100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011110001000011101100111011101110110011001100100010101010101010101010100001100110011001100110011001000100010001000100010000100010010000100100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000100010001100110011010001000100010001000101010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111011101100110011001100110011001100110011001100110011001100110011001100101010100110011001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000110011001100110011001100110011010001000100010001000100,
	2400'b010001000100010000110010000100100001000100010001000100010001001000010001000100100011001000100010001000110011001000110011001101000100010001000100001000010001000100010001001000100010001001010110011101110110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100100001100100010001000100010001000100010001000100010001000110011010001100101011001100110011001100110011101110111011101110111011101110111011101100100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001110111011101110111011001110110011101110111011101110111011101110111011001100110011001000100010001000101011001010110011001000100001100110100001100110100001100110011001100110011001101000101010001010100010001000100010101100110011001100110011001100110011001100110011101100110011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100110011001100110010101010110011001100111011101110111011001110111011001100111011001010101010101100110010101010100010000110011001100110010001000100010001000100010001000010001001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000100011010001000100010001000100010101010101011001100110011001100110011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110110011101100110011101100110011001100110011001100110011001100110011001100110010101000011001000100010001000100010001000100010001000100010000100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001100110011001100110011010001000011010001000100010001000100,
	2400'b010101000100001100100001000100010001000100010001000100010001001000010001001000100011001000110010001000110011001100110011001100110100010001000011001000010001000100010001000100100010001001100111011101110110011101110111011101110111011101110111011101110111011101110111011101100111011001100110011001100100001100110010001000100010001000100010001000100010001000100011010001010110010101100110011001100110011101110111011101110111011101110111011101110101010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101100110011101110111011101110111011101110111011101100110010001000100010001010101011001100110010101000100001101000011001100110100010000110011001100110011001100110100010101010100010101010100010101100110011001100110011001110110011001100110011001100111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100110010101010101010001000100010001000101010101100101010101100101011001010101001100110011010001000100010001000100010000110011001100110010001000100010001000010010001000100001001000010001001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001100110100010001000101010001000100010101010110011001010110011001100110011001100110011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101100110011001100110011001100110011001100110011001010011001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001100110011001100110011010001000100010001000100010001000100,
	2400'b010001000100001000100001000100010001000100010001000100010010001000010001001000110011001100110010001101000100001100110100001100110100010101000011000100010001000100010001000100010001001101100110011001110110011101100111011101110111011101110111011101110111011101110111011101110111011001100110011001100100001101000011001000100010001000100010001000100010001000100011010001010110011001100110011001010110011001110111011101110111011101110111011101110110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110110011101110111011101110111011101100111011001100100010001000100010001010110011001100110010101000100010001000100001101000100010000110011001100110011001100110100010101010101011001100101010101010110011001100110011001100110011001110111011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100110010101010101010101000100010001000100010000110011001101000100010001000011001100110011001000100010001000100011010001000100001100110011001000100010001000100010001000100010001000010001001000100010000100010010001000100010001000100010001000100010001000100010001000100010001000100011001101000100001101000100010001010101010101010101010101100110011001010100010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101100111011001100110011001100110011001100110011001100100001100100010001000100010001000100010001000100010001000100010001000100010001000010010000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000110011001101000100010001000100010001000100010001000100,
	2400'b010001000011001000100001000100010001000100010001000100010010001000010001001000110100001100110011001101000100010000110100010000110100010001000010000100010001000100010001001000010010010101110110011001110111011101110110011101110111011101110111011101110111011101110111011101100110011001100110011001100100010101010011001000100010001000100010001000100010001000100010001101000101011001100110011001100110011001110111011101110111011101110110011101110110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011001010100010001000100010001100110011001100110010001000100010001000100010001000100010000110011010000110011001101000100010101010101010101100101010001010101011001100110011001100110011101110110011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110110011101100110011001010101010101010101010001000100010001000100010001000100001101000011001100100011001100100010001000100010001000110011001100110010001000100010001100100010001000010001001000100001000100100010001000010001000100010010001000100010001000100010001000100010001000100010001000110011001100110100010001010101011001100110010101010110010101010101010001000101010101010110011001100110011001100110011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110010101000010001000100010001000100010001100100010001000100010001000100010001000100010001000100001000100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100011001101000100010001000100010001000100010001000100,
	2400'b010000110010000100010001000100010001000100010001000100100010000100100010001000110100001100110011001101000101010000110100010000110011010101000010001000010001000100010001000100100011011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101010110011101100110011001010100011001010100001000100010001000100010001000100010001000100010001000110101011001100110011001100110011001100111011101110111011101110111011101110110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011001100110011001000100010001000101010101100111011101100101010001000100010101000100010001000100010000110100010101000011001100110100010101010101010101100110010101010101011001100110011001100110011001110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001100111011101100110011001100110011001010101010101000100010001010100010101000100010001000011001100110011001100100010001000100010001000100010001100110011001000100010001100110010001000100010001000100010001000100010001000100010000100100001001000100011001000100010001000100010001000100010001000100011010001000101011001100101010101000101010001000100010000110011001101000100010001000101010101010101010101100110011001100110011001100111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001101000100010001000100010001000100010001000100,
	2400'b010000100001000100010001000100010001000100010001000100100010001000100011001101000100010000110011001101000101010100110100010001000011010101000010001000010001000100010001000100100100011001100110011001100110011101110111011101110111011101110111011101110111011101110111011001010111011101100110011001010101011001100100001000100010001000100010001000100010001100100010001000110011010101100110011001100110011001100111011101110111011101110111011101110110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110110010001000100010001010101010101100111011101010101010001000100010101010100010001000100010000110100010101000100010001000100010101100101010101100111011001010101010101100110011001100110011001110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011001110111011001100110011001100110011001100101010101010100010001010101011001010101011001010100010001010100001100110011001100110010001000100010001000100011001100110011001100110011001100100010000100100010001000100001001000100010000100010010001000100010000100100010001000010010001000100010001101000101010101010101010101000011001100110011001100100010001000100010001100110011001100110100010001000100010001010101010101010110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110010101000010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000110100010001000101010101000101010101010101,
	2400'b001000100010000100010001000100010001000100010001001000100010001000100011001101000100010000110100001101000101010101000100010001000011010001000010000100010001000100010001000100100101011101100110011001100110011001110110011101110111011101110111011101110111011101110111011001110111011101110111011001010110011001100100001100110010001000100010001000100010001100100010001000100011010101100110011001100110011001100111011001110111011101110111011101100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101100101010001000101010101010101011001100111011001010101010001000101010101100100010001000100010001000101010101010100010001000100010101100101010101100111011101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101100110011101110111011001100101010101010101010101010110011001010110011001010100010001000011001100110011001101000100001100100010001000100010001000110011001100110100001100110010001000010010000100100001000100010001000100010010001000100010001000100010001000100010001000110100010001010101010101000011001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001000100010101010101011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100101010000100010001000100011001000100010001000100010001000100010001000100010001000100010001000110011001100100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100011010001000101010101010101010101010101,
	2400'b001000100001000100100001000100010001000100100010001000100010001100100100001101000101010000110100001101000101010101010100010001010100010001000010000100010001000100100001000100110110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110110010101100110011001100100010000110010001000100010001000100010001000100010001000100011010001010110011001100110011001010110011101110111011101110111011101100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011001010100010101010101010101010110011001100111011001100101010001010101011001100101010001000100010001000110011001010100010101000101010101100110010101010110011101100101010101100110011001100110011001100110011001110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010110011001010110011001100111011101100101010101000100010001000011010001000011010001000011001100110011001000100010001000100010010001010100010001000100001100100010001000110010001000100001000100010010001000100010001000100010001000100011001101000100010001000011001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110100010001000100010101010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011001100110011001100110011001100100001000100011001000100010001000100010001000100010001000100010001000110011001100110011010001000011001100100010001000100010000100100001000100010001000100010001000100010001000100010001000100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001001000101010101010101010101010101,
	2400'b001000010010001000010001000100010001000100010010001000100010001100110100001101000101010101000100010001000101011001010100010101010101010001000010000100010001000100100010001001000110011001100110011001100110011001100110011001110111011101110111011101100111011101110111011101110111011001100110010101100110011001100100010000110011001000100010001000100010001000110010001000100011001101010110011001100110011001100110011101110111011101110111011101110110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001110111010101000101010101010110011001100110011101100110011001100101010001010101011001100101010001000100010001010110011001100100010101000101010101100110010101010110011001110110010101010110011001100110011001100110011001100110011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001010110011001100101010101100101010101010101010101000100010001000011001100110100001100110010001000010001001001000101010101010101010101000010000101000100001000100010000100010001000100010010001000100010001000110011001101000011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011010001000101010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001000010001000110011001000100010001000100010001000100010001000100011001100110100010001000100010001000100001100100010001100100010001000100010001000100010000100010001000100100010000100100010001000100001000100010001000100010010001000100001000100010001000100010001000100010001000100010001000100010001000100010001001000100011010001010101010101010101,
	2400'b001000100010000100010001000100010001000100100010001000100011010000110100001101000101010101000100010001000101011001100101010101010101010100110010001000010001000100010010001101100110011001100110011001100110011101110111011101110111011101110111011001100111011101110111011101110111011101100101011001100110011001010100010101000100001000100010001000100010001000100011001000100010001100110101011001100110011001100110011101110111011101110111011101110110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110110011001100110010101010110011001100110011001100110011001100110011001100101010001010101011001110110010001000100010001100111011101100101010101000101011001100110011001010110011001100110010101010110011001100110011001100110011001100110011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011001110110011001100110011001100110011001010101010101010100010001000100010001000011001100110011001100110100001101000011001100100010001000100011010101010110011001010011000100110110001101000100001000100001000100010010001000010010001000100010001000100010000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010001010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110010000100010001100110011001000100010001000100010001000100010001000110011001101000100010101010100010101010100001100100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001100100010001000100010000100010001000100010001000100010001000100010001000100010001000100010010001101000100010101010101,
	2400'b001000100001000100010010001000010001001000100011001000100011010000110100001101000101010101010100010001000101011001100110010101010101010100110010000100100010000100100010010001100110011001100110011001110111011101110111011101110110011001110111011001100110011001110111011101100110011101100110011001100110011001010101010101000100001100100010001000100010001000110010001100100010001000110100011001100110011001100110011101110111011101110111011101110110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100101011001100110011001100110011001100110011001100110011001100101010001100110011001110110010101000101011001110111011101100101010101010101011001100111011001010110011001100110011001010110011001100110011001100110011001100110011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100110011001100110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110110011001100110010101010100010000110011001100110011001100110011001100110010001100110011001100110100001100110100010001000011001000010001001101010110011001010101001000100101001001000100010001000010000100010010000100010010001000100010000100100001000100100010000100100001001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001000101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100100001100110011001100100010001000100010001000100010001000100011001100110100010001000101010001010101010101010100010000110010001000100001000100100011001000010001000100010001000100010001000100010001000100010001000100010001000100010010001100100010001000110010001000100010001000010001000100010001000100010001000100010001000100010001000100100010010001010101,
	2400'b001000100010001000100010000100010010001000100011001000100100010000110100001100110101010101010101010001010101011001100110011001100101010101000010000100100010001000100011011001110110011001100110011001110111011101110111011101110111011101110111011001100110011001100110011001110110011001100110011001100110011001010110010101010101001100100010001000100011001000110010001100110010001000110100010101100110011001100110011101110111011101110111011101110110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110010101100110011101110110010101000110011101110111011101110101010101010101011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001110110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100111011101100110011001100110011001100111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100001100110011001100110011001100110011001100110011001100110011001100110011001100110100001100110011001100110100010000110010000100100100011001100101001100010011001001000100010000110010001000100010000100010001001000100001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110100010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001000011001100110011001100100010001000100010001000100010001000110100010000110101010101000101010101010100010001000100001100110010001000100010000100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001100100011001100110011001100100010000100100010000100010001000100010001000100010001000100010001000100010010001001000101,
	2400'b001000100010001000100010001000100010001000110011001000110100010000110100001100110101011001100101010001010101011001100110011001100110010101000010000100010010001000100011011001110110011001100110011001110111011101110111011101110111011101110110011001100110011001110110011001100110011001100111011101100111011001010110011001100101001100100010001000100010001000110011001000110011001000110011010001100110011001100110011101110111011101110111011101100111011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110010101100110011101110110010101010111011101110111011101110110010101010110011001100111011101100110011001100111011001100110011001100110011001100110011001100110011001100111011101110111011001100110011001100110011001100110011101100110011001100111011001100111011001100111011101100111011101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010000110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010000110011001101000011001000010010010001010101001100010010001000110100001000010010001000100001000100010001000100100001000100010010001000010001000100100010001000100010001000100010001100110010001000100010001000100010001000100010001100110011001100110011001100110011010001010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010000110011001100110011001000100010001000100011001000110011001100110101010101010101010101010101010101010101010101010011001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100110011001100110011001100010001000100100010000100010001000100010001000100010001000100010001000100010010001000100011,
	2400'b001000100010001000100010001000100010001100110011001000110100010000110101010000110101011001100101010101010110011001100110011001100110011001010010000100010001001000100100011101110110011001110110011001110111011101110111011101110110011001100111011001100110011001100110011001100110011001110111011101110110010101100110011001100110010000100010001000100010001000110011001000100011001100110011001101000110011001100110011101100110011001110111011101100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011101100110011001100110011001010110011001100110011001100110011001100110011101110110010101100111011101110111011101110101010101010110011001100110011001100110011001100110011001100110011001100111011001100110011001100110011001100111011101110111011101100110011001100111011101100110011101110110011001100110011001100110011001100110011101110111011001100110011001110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000100010001000100010000110100001101000011010001000011001101000100010101010101010101100110011001100101010101010101010101010100010000110010001100100001000100110100001100010001000100100010000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000110011001101000100001100110011001100110011001000110011001100100011001100110011001100110011001100110101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100100001100110011001100110011001000100010001000100011001100110011001100110101011001100110010101010110011001010101010101010100001100100010001000010001001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010010000110011001100110010000100010001001000100001001000100001000100010001000100010001000100010001000100010001000100010010,
	2400'b001000100010001000100010001000100011010000110011001000110101010000110101010000110100011001100110010101010110011001100110011001100110011001100011000100010001001000100101011101110111011001100111011101110111011101110111011101100111011101100110011001110111011001100110011001110110011001110111011101110110011001100110011001100110010000110010001000100010001000110011001000100010001100110011001101000101011001100110011101110110011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110011101110110011001110111011001100110011001100110011001100110011001100110011101110110010101100111011101110111011101100110011001010110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011001100110011001100111011001100110011001110111100010001000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010001000100010001000100010001000100010001000100010101000100010001010101011001100110011001100110011001010101010101010101010101000101010101010101010000110010000100010010001000100001000100010001001001000011000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000110011001101000100010001000100010001000100001100110100001100110010001000110011001100110011001100110100010101100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001000011001100110011001100100010001000100010001000110011001100110011010000110100011001100110011001100101011001010101010001000100001100110010001000010001001100100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010010001000011001100100001001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010010,
	2400'b001000100010001000100010001000100011010000110011001100110101010001000101010100110100011001100110011001100110011001100110011001100110011001100101001000010001001000110110011101100111011001110110011101110111011101110111011101110111011101100110011001100110011001100110011101100111011101110111011101100110011001100110011001100110010001000011001000100010001100110011001000100010001100110100010001000100011001100111011001110110011101110110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101100110011101110111011001100110011001100110011001100110011001100110011001110110011001110111011101110111011101100110011001100110011001100110011101100110011101100110011001100110011001100110011001100110011101100110011001110111011101110111011101100111011001100111011101110111011101110111011101110111011101100111011101110111011101100110011001100111011101111000100010001000011110001000100001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000100010001000100010001000100010001010101010101010101010101010101010101010110011001110110011001010101011001010101010101000100010001000011001101000100010101010011000100010001000100010001000100010010010101100011000100010001000100010001000100010001000100010001000100010010001000100010001000110010001000100011010001000100010001000100010101000100010101000100010001000011001000110011001100110011001100110011010001010111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110010100110011001100110011001000100010001000100010001000110011001100110011010001000100010001100111011001100110011001010101010001000011001100100010001000100010001000010001001000010001000100010001000100010001000100010001000100010001000100010001000100010010010001000011001000100010001000100010001000100010001000100010000100010001001000010001000100010001000100010001000100010010,
	2400'b001000100010001000100010001000110100001100110011001100110100010001000101011001000011010101100110011001100110011001100110011001100110011001100100001000100010001000110110011101100111011001110111011001110111011101110111011101110111011101100110011001100110011001110111011001100111011001010110011101100110011001110110011101100110010101010011001000100010001000110011001100100010001100110100010001000100010101100110011101100110011001100110011001110111011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101100111011101110111011001110111011101110111011001100110011001100110011001100110011001100110011001100101011001110111011101110111011101110110011001100110011001110111011101110111011001100110011001100110011001100111011001110111011101100111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101100110011001100110011001110111011110001000100010001000011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010100010001000101010101010101010101010101010101010110011001010110011001100110011001110110011001000100010000110011001100110010001000100010000100100010001000110100001100100001000100010001000100010011011001010010001000100001000100010001000100010001000100010001000100010010001000100010001000110011001100110011010001010101010101010101010101010100010101100101010101010100001100110101010000110011001101000100010001000110011101110111011101110111011101110111011101110111011001110111011101110111011101110111011001100101001100110011001100110011001000100010001000100010001100110011001100110100010001010101010101010110011101100110011001010100010001000011001100110010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100100100010001000011001101000011001100110011001100110010001100100010001000100010001000010001000100010001000100010001000100010001,
	2400'b001000100010001000100010001001000101001100110011001101000100010001010101011001010011010101100110011001100110011001100110011001100110011001100100001000100010001001000111011101100111011101110111011101110111011101110111011101110110011101100110011001100110011001110111011001100111011101100110011001100111011101110110011001100110010101010100001100100010001000110100001100100011001100110011010001000100010101100110011101110111011101100111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100101011001100111011101110111011101110110011001110111011001110110011001110111011001100110011001100110011101110111011101110111011101100111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110110011101110110011001100110011001110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110110010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110010101010100010000110011001000100010001000100010001000010001000100010001000100010010001101000010000100010001000100010010001100100001001000100010000100100001000100100010001000010001000100010010000100100010001000100010001100100011010101100101011001100110011001100101010101100110011001100110010101010110011001010100001101010110010101000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001010011001100110011001100110010001000100010001000100011001100110100010001000100010001010110011001100110011001100110010101010101010001000100001100110010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100100100010001000101010001000100010001000100001100110011001100100011001000100010001000010001000100010001000100010001000100010001,
	2400'b001000110010001000100010001101000100001101000011001101010100010001010101011001100100010101100110011001100110011001100110011001100110011001100011000100100010001001010111011101100111011101100110011101110111011101110111011101110111011101100111011101110111011101100111011101110111011101110110011001110111011101100110011001100110010101010100001100100010001000100011010000110011001100110011010001000100010001100110011001110111011101100111011101110110011001100110011001100110011101100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101100111011101110111011101110111011101110111011101110110010101100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101011001010110011001100110011001100110011001100110010101010110010101010101010000110011001000100010001000100010001000100010001000010001000100010001000100010001000100100011001000010001000100010001000100010010010000110011001000110010001000100010001000100010001000010001000100010010001000100010001000100011010001010101010101100110011001100110010101100110011001100110011001100110011001100110010101010110011101100101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001100100010001000100010001100110011010000110100010001000101010101010110011001100110011001100110010101010101010101000100001100110010001000110010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010101000100010001000100010101000100010000110011001100110011001000110011001000100010000100010001000100010001000100010001,
	2400'b001100110010001000100010001101010100001100110011010001010100010001010101011001100101010001100110011001100110011001100110011001100110011001100011000100100010001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001110111011101110111011101110111011101110111011101110111011001100110011001010100001100100010001000100011010000110011001100110011010001000100010001010110011001110111011101110110011001110111011001100110011001100110011001100111011101100110011101100110011001100110011001100110011001100111011101100110011101100110011001100111011101110111011101100110011001110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010000111100010001000100001110111011101110111011101110111011101110111011101110111011101010101010101100110010101100110011001100110011001100110011001100110011001100101010101010101010000110011001100110011001000100010001000100001000100100010001000010001000100010001000100010001000100010010000100010001000100010001000100100011010001010100010000110011001100100011001100110011001000100010001000100010001000100010001000100010001000110011010001010101010101100110011001100110011001100110011001100110011001100110011001100110011101110110010101010110011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110011001000100010001000100011001100110011010001000100010101000101011001100110011001100110011001100110010101010101010101010101001100100010001000110010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010101010101010101010101010101010101010001000011001101000011001101000011001100110010001000010001000100010001000100010001,
	2400'b001100110010001000100010010001010011010000110100010001010100010001100101011001100110010001100110011001100110011001100110011001100110011001100010000100100010001101100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011001100110011001010100010000110010001000110011010000110010001100110100010001000101010001000110011001110111011001110111011101100110011001100110011001100110011101110110011001100111011001100110011001110110011001100110011001100111011101100110011001110111011101100110011001110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000100010000111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100101010101010100010001000011001100110011001100110011001100110010001000100010001000100001000100010010001000100001000100100010000100010001000100010001000100010001000100010001000100010010001101000101010000110011001000100010001000100010001100100011001100100010001000100010001000100010001000100010001100110011010001000100010101100110011001100110011001100110011001110111011001110111011001110111011001010101011001110111011101110111011101110111011101110111011101110111011101100100001100110011001100110011001000100010001000110011010001000011010001000100010101010101011001100110011101110110011001100110010101010101010101010101010000100010001100110010000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100100010101010101010101010101010101010101010101000100010001000011010001000011001100110011001000100010001000100001000100010001,
	2400'b001100110010001000100011010001010011010000110100010101010100010001010101011001100110010101100110011001100110011001100110011001100110011001010010001000100010010001100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001100110011001100110011001100101010000110011001100110100010000110010001100110100010001000101010001000110011101110110011001110111011001100110011001100110011101110111011101110110011001100111011001100111011001110111011101100110011101100111011001110111011101110111011101110110011001100110011001110111011101110111011101100110011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110110011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110010101010100010000110011010000110011001100110011001100110011001100100011001000100010001000100001000100100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100100010001000100010000100010001001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100011010001000101010101100110011001100110011001100111011001110111011101110111011101100110011001100111011101110111011101110111011101110111011101110111011101000011001100110011001000110010001000100010001101000011010001000100010001000101011001100110011001100111011101100110010101010101010101010101010101010101010000100010010000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010100010101010110011001100110010101010101010001000100010101000100010101010100010001000011001000100010001000100001000100010001,
	2400'b001100110010001000100011010101010011010000110100010101100100010001010110011001110110011001010110011001100110011001100110011001100110011001000001001000100010010101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001110110011001100110011001100110011001100101010100110011001100110100010001000011001101000100010001000101010101000101011001100110011001110110011101100111011101100110011101110111011001110111011101100110011001100110011001100110011001110111011101110111011101110111011101110111011001110111011001110110011101110111011101110111011001100110011101110111011101100101011001100110011001100110011001100110011001100110011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001010101010001000011001101000100010001000100010000110011001100110011001100110011001000100010001000100010001000100010001000010001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100001000100100010001000010001000100100010001000100010001000100010001000100010001000100010001000100010001000110011010001000101011001100110011001100110011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111010100110011001100110011001100110010001000110011001101000100010101010100010001010101011001100110011001100110011001100101010101010101010101010101010101010100001100100010001100110011001100100001000100010001000100010001000100010001000100010001000100010001000100010010000100100010010001010110010101010101010101010101010101010101010101000101010101010101010001000100001100100010001000100001000100010001,
	2400'b010000110010001000100011010101010011010001000100011001100100010101100101011001110111011001100110011001100110011001100110011001100110011000110001001000100011010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110010101000011001100110100010001000011001101000101010001000100010101000100011001100111011101110110011101110111011101110110011001110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101100111011101110111011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100101010001000100010001000011010001000100010001010100010000110011001100110011001100110010001000100010001000100010001000100010001000010010001000100001000100010001000100010001000100010001000100010001000100010001000100100010010001000100001100110010000100100010001000010001000100010001000100010010001000100010001100100010001000100010001000100010001000110010001100110011010101100110011001100111011101110111011101110111011101110110011101110110011001110111011101110111011101110111011101110110001100110011001100110011001100110011001000110011010001000101010101000101010101100110011001100110011001100110011001100110011001100110011001100110011001100100001000100010010001000011001100100010000100010001000100010001000100010001000100010001000100010001001000100010001000100010001101000101010101100110011001100101010101010101010001010101010101010101010001000100001100110010001000100010001000010001,
	2400'b001100100010001000110100010101010100010101000100011001100100010101100110011001110111011101100110011001100110011001100110011001100110011000100001001000100011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110010101000011010001000100010001000011001100110101010101010101010101000100011001100110011101110111011001110111011001100111011001110111011101110110011101110111011101100110011001110111011101110110011001110111011101110111011101110111011101110111011101110111011101100111011101110111011101100101011101110111011101100110011001100110011001100110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110010101010100010001000100001100110100010001010101010101010100001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100100110011001100110010101000010001000100001001000010001001000010001000100010001001000100010001100110011001000100010001000100010001100110010001000100011001101000110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100100011001100110011001000110011001101000100010101010100010101010101010101100110011001100111011001100110011001100110011001100110011001100110011001100101001100100011010101000011001100110010000100010001000100010001000100010001000100010010001000100010001000100010001000100011010001000101010101100110011001100110010101010101011001100101010101010100010001010100010000110011001100100010001000100001,
	2400'b001100110010001000110100010101010101010101010101011001100100011001100110011001110111011101100110011001100110011001100110011001100110010100010001001000100100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000011001100110100011001100110010101000100010101100110011001110111011001110111011001100111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101011001110111011001100101011001110111011001010110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011001100101010101010100010001000100010001000100010101010101010101000010001100100010001100110011001100100010001000100010001000100010001000100011001000100011001000100010000100010001000100010001000100010001000100010001000100100010001000100100011101110111011001000010001000100010001000100010001000100001000100010010001000010001001000100011001000110011001000100010001100110010001000100011001100110100011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001100110011001100110011001101000100010101010101010101010101011001100110011001110111011101110110011001100110011001100110011001100110011001100101001000100100010101000010001100100001000100010001001000100001000100010001000100010001001000100010001000100010001000100010010001010101010101100110011001100110011001100110011001100110010101010100010101010100010000110011001100100011001000100001,
	2400'b001100110010001100110100011001010101011001010101011001100100010101100110011001110110011101100110011001100110011001100110011001100110010000010001000100100101011101100111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101000100010001010011001100110100010101100110011001010100010101100110011001110110011101110111011101110111011101110111011101110111011101110110011001110111011101100111011101110111011001110111011101110111011101110111011101110111011101110110011001100101010101110111011101110101011001110111011001010110011001100110011001100110011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010000111011101110111100010001000100001110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011001100101010101010101010001010100010001000100010101010101010000110011001100100010001100110011001000100010001000100010001000100010001100110011001100100011001000100001000100010001000100010001000100010001000100010001000100100010001000100010011010001000011001000011001000110010001000100010001000100010000100100010001000010001000100010010001000100010001100110011001100110010001000100011001100110011010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001100110011001100110011001100110011010001000100010101010101010101100110011001110111011101110111011101110111011101100110011001100110011001100110011001100101001000100101010100110010001000010001000100010001001000100001000100010001000100010001000100100010001000100010001000100010001101000101011001100110011001100110011001100110011001100110010101010101010101010101010001000011001100110011001000100010,
	2400'b001100110011001101000100011001100101011001100101011001100101011001100110011001100110011101100110011001100110011001100110011001100110001100010001000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000100010001010011001100110011010101100110011001100110010101100110011001100111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101010110011101110101010101100111011001100110011001100110011001100111011001100110011001100110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101111000100001111000100010000111100001110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101010101010001010101010101010100001100110011001100110011001100110010001000100010001000110010001000100011001000110100001100110010001000100001000100010001000100010001000100010001000100010001000100100011001000100010001001101000011001000011001000110010001100110010001000100010001000100010000100010010001000100010000100010010001000100011001100110010001000110010001100110011001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110011001100110011001100110011010001000101010101010101010101100110011001110111011101110111011101110111011101100110011001110111011001100110011001100100001000100101010000100010001000010001000100010001000100010001000100010001000100100010000100100010001000100010001000100011001100110100010101100110011001100110011001100110011001100101010101100110011001010101010101000100010000110011001100110010,
	2400'b001100110011001101000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000010001000100110110011001100111011101110111011101110111011101110111011101110111011101110111011101110110011101110110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000101010001000011001100110011010101100111011101110110010101100111011001100111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001110101010101100110010101100110010101100110011001100111011001100110011001100110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000011110000111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100101010101010100010101010101010100110011001100100011001100110010001000110011001000110010001100110011001000110011001100110100010000100010001000010001000100010001000100010001000100010001000100010001000100010010001100110011001000100110011101000010001100110011001100110011001000100011001100100010001000100010001000100001001000010010001000100010001100110011001100110011001100110011001100110101011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110011001100110011001100110011001101000100010101000101010101100110011001100110011001110111011101110111011101110111011101100110011001100110011001100110011001100100001000110101001100100010000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000110011010001010101010101010101011001100110011001100110011001100110011001100110011001100101010101000101010001000100001100110010,
	2400'b001100110011001101000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001000101000110011001100111011101110111011101110111011101110111011101110111011101100110011101110111011101100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101000011001100110011010001100111011101100111011001100110011001100110011001110111011101100111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101100110011001100101010001100101010101100101010101010101011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101100110011001100110010100110100010101010100001100110011001000100011001100110010001000110011001100110011001100110011001100100100001100110011001000100010001000100001000100100001000100010001000100010001000100010001000100010001001000110011001100100010011001010100001101000011010001000011001101000011001100100011001100100010001000100010001000100001001000100010001000100011001100110011001100110011001100110011010101110111011101110111011101110111011101110111011101110111011101110111011101100011001100110011001100110011001100110011010001000100010101010110011001100110011001100111011101110111011101110111011101110111011101110111011101100110011001100110011001100100001000110101001100100010000100010001000100010001000100010001000100010001000100100001001000100010001000100010001000100011010001010101010101100110011001100110011001100110011001100110011001100101010101010101010101010101010001000100001100110010,
	2400'b010000110011001101000101011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100011000100010001000101000111011001100111011101110111011101110111011101110111011101110111011101100110011101110110011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001010101010101000011001100110011010001100111011101100111011001100110011001110111011001110111011101110111011101110111011001110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010110011001010101010001010101010101010101010101010101011001100110011001100111011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101111000100010001000100010001000100010001000100010001000011101110111011101110111100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100101001100100011010001000011001100110011001000110011001100110011001000110011001100110011001100110100010000100011001100100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001001000110011001100110010001001010101010101010100010001000011010001000100001100110100001100110010001000100010001000100010001000100010001000100010001101000011001100110011001100110011001101010110011101110111011101110111011101110111011101110111011101110111011101000011010000110011001100110011001100110100010001000101010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011001100110011001100011001001000100001000100010000100010001000100010001000100100001000100010001000100100010001000100010001000100010001000110011001101000101010101100110011001100110011001100110011001100110011001010101010101010110011001010101010001010100010000110011,
	2400'b010001000011010001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000100010001001001010111011001100111011001110111011101100111011101100110011101100110011101110111011001100110011101110111011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001010110010101000100001100110011010001100111011001100111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101001101000100010101010100010001010101011001100111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001010011001000100010001100110011001100110011001100110011001100110100001100110100010001000011010001000100010000110011001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100100011001100110011001000110101011001100101010101000100010001010100001101000011010000110011001100110011001000100010001000100010001000100010001000110011001100110011001100110011001100110100011001110111011101110111011101110111011101110111011101110111011000110011010000110011001100110011001101000100010001010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011001100110011001100011001000110011001000100010001000010001000100010001001000100001000100010001000100100010001000100010001000100010001100110100010001000101010101100110011001100110011001100110011001100110011001100110011001100110011001010101010101010100010000110011,
	2400'b010001000100010001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010001000100010001001001010111011001100110011001100110011001100111011001100110011001100110011101110111011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110010101000100001100110011010001100111011001110111011001100110011001100110011001100110011101110110011001100111011001100110011001100110011001100110011001100110011001100110011001100111011101100111011101110111011101110111011101110111011101100110011001010100010001010100001100110100010101000101010001010110011001100110011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011101100110010100110010001000100011001100110011001100110011001100110011001100110100001101000100010101010100010001000011001100100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001100110011001100100010010101100101011001010101010101000100010001000011010000110011001100110011001000100010001000100010001000100010001000100011010001000011001100110011001100110011010101100111011101110111011101110111011101110111011101110110010000110011001100110011001100110011001101000101010101010110011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001100011001000110011001000100010000100010010000100010001001000100001000100010001001000100010001000100010001000110011001100110011010001010110011001100110011001100111011101110110011001100110011001100110011001100110011001100101010101010101001100110100,
	2400'b010001000100010001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000001000100010001001101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001100110010101000100001100110011010001100111011101100111011001100111011101110111011101110111011101110110011001100110011101110110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110110011101100110011001010100010101000100001100110100010001000100010101010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011001100101001100100010001000100011001100110011001100110011001100110011001100110100010001010100010001010101010101010100001100100010001000100011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000110011001100110010001101100110010101010101010101010100010001000100010000110011010000110011001100110010001000100010001000100010001000100010001101000100001100110011001100110011010001010110011101110111011101110111011101110111011101110101001100110011001100110011001100110011010001010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100011001000110010001000100010000100100010001000100010001000100010000100010001001000100010001000100010001000110011001101000100010101100110011001100110011001110111011101110110011001100110011001100110011001100110011001010101010101010101001101000100,
	2400'b010101010100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001000100010010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110010101000101001100110011010001010111011101100111011001100111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011101110110011001110111011101110111011101110111011001100110011001100101010101010100001100110011001100110100010001010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100011001000100010001000110011001100110011001100110011001100110011001100110100010101010110011001010101010101010100001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011010000110010001001000110011001100110010101010101010101000100010001000100010001000011001100110011001000110011001000100010001000100010001000100011010000110011001101000100010000110100011001110111011101110111011101110111011101100100001101000011001100110011001101000100010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011001010011001100110010001000100001001000100010001000100010001000100010000100010001000100100010001000100010001100110011010001000101010101100110011001100110011001110111011101100111011101100110011001100110011001100110011001010101010101010100010001000100,
	2400'b010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100001000100010010010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101001100110011010001010110011101110111011001100111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011101110110011001100110011001100110011001100101010001000101001100100011001000110011001101000101011001100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010100110010001000100010001000110011001100110011001100110011001100110011001101000101010101100110011001100110010101010010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010010001000011001000100101011001100110011001100101010101010101010001000100010001000100001100110011001100110011001000100010001000100010001000100010001101000011001101000100010001000011010101100111011101110111011101110111011101010011001101000011001100110011001101000100010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010011001100110010001000100010001000100010001000100010001000110010000100010010001000100010001000100010001100110011010001000100010101010110011001100110011101110110011101100111011101100110011001100110011001100110010101010110010101010100010001010101,
	2400'b010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000010001000100010010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010000110100010001100110011101110111011001100111011001110111011101110111011101110110011001100111011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110110011001100111011001100110011001100101010101010100010000110100001100100010001000110011001101000100011001110110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101001100100010001000100010001100110011001100110011001100110011010000110100010001010101011001100110011001100110010000110010001000100010001000010001000100010001000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001001001000100001000100011011001100110011001010110010101010101010101010100010001010100010000110100001100110011001100110010001000100010001000100010001000110011001100110100010001000100010001010110011101110110011001100111011001010011010001000011010000110011010001000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011001010010001100100010001000100010001000100010001000100010001100110010000100010010001000100010001000100010001100110011001101010100010101100110011001100110011101110111011101110111011101110110011001100110011001100101011001100110011001010100010101010101,
	2400'b010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110001100010001000100010011011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110010001000101010101100110011001110111011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011001100110011001100110010101010100010101000100001100110011001100100010001000100011001100110101011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010011001000100010001000100010001100110011001100110011001100110011010001000100010101010101011001100110011001110101001100100010001000100010001000010001001000010001000100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100100100001100100010010001100111011001100110011001100101010101010101010101010101010001000011001100110011001100110011001000100010001000100010001000110011001100110100010001000100010001000101011001100110011001100110011001000011010001000100010001000100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011001000010001100100010001000100010001000100010001000110010001100110010000100010010001000100010001000100011001100110011001101010101010101100110011001100110011101110111011101100111011101110110011001100110011001100110011001100110010101000101010101010101,
	2400'b010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100101001000010001000100100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000101010101100110011001110111011101110111011101110111011101110111011101100110011101110111011101100110011001100110011101110111011101110110011101110111011101100110011001110111011001100110011001100110011001100110011001010100010001000100001100110011001100100010001000100011001100110101011001010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010100110010001000100010001000110011010000110011001100110100001101000100010001010101010101100110011001100101010101000011001100100010001000100010001000010001001000010010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100100010001101010111011101110110011001100101011001100101010101010101010101000100001100110011001100110011001000100010001000100010001000110011001100110011010001000100010001000100010101100110011001100110010101000100010101000100010001010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001000011001100100010001000100010001000100010001000100011010001000011000100100010001000100011001000100011001100110100001101000110011001010110011001100110011001110111011101110111011101110110011001100110011001100110011001100101010001010101010101010101,
	2400'b010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001001000100101011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100111011101110111011001100110011001100110011101110111011001100110011001100110011001100110011001100110011001100110011001100110010101000101011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101100110011001100110010101010100010000110011001100110011001100110010001000100011001101000101010101000101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100100010001000100010001000110100010001000100010001000100010001010101010101010101011001100110011001100110010101000011001100100010001000100010001000010010001000100010001000100010001000010001000100010001000100010001000100100001000100010001000100100010001000010001000100010010001100110010001001000111011101110110011001100110011001100110011001100101010101010101010000110100010000110011001100100010001000100010001000110011001101000100010001000100010001000100010101010110011001100110010100110100010101000100010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001000100010001000100010001000100010001100110011010000110010001000100010001000100011001100110011001101000100010001000110011001100110011001100111011101110111011101110111011101110110011001100110011001100110011001010101010101100101010101010101,
	2400'b010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100011000100010001001000110110011001100110011001100110011101100110011101100110011001100110011001100110011001100110011001100111011001110111011001110111011001100110011001100111011001110111011101100110011001100111011001100110011001100110011001100110011001100110010101000101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010101100110011001100110011001100110010101000101010000110011001100110011001100100010001000100011001101000100010001010110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011001010011001000100010001000100010001100110101010001000100010001000101010101010101011001100101011001100110011001010101010000110011001100100010001000100010000100010010001000100010001100100010001000010001000100010001000100010001001000100001000100010001000100100010000100100010001000010001001000100010001000110110011101110111011101100110011101100110011001100101010101010101010101000100010001000011001100110010001000100010001100110011001101000100010001000100010001000100010101010101011001100110010000110100010101000101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110011001000100010001000100010001000100010001100110011010000110010001000100010001000100011001100110011001101000100010001000110011001100110011001110111011101110111011101110111011101110111011101100110011001100110011001010110011001100101010101010101,
	2400'b010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010010000100010001001000110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011001110111011101110111011001100110011001100110011001100111011101110111011001100110011101100110011001100110011001110110011001100110010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001010101010001000100010001000100010001010110011001010101010001000011001100110011001100110011001100110010001000100011001100110100010001010101011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110010001000100010001000100011001101000101010001000100010001010110010101100110011001100110011001110111011001000100010000110100001100100010000100010010001000100010001000100011001100110010001000010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000110101011001110111011101100110011101100110011001010101011001010101010101010101010001010100001100110010001000100010001100110011001101000100010001000100010001000100010001010101011001100110010001000101010101010110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001000100010001000100010001000100011001100110011001100110010001000010010001000100011001100110011010001000100010001000110011001100110011001110111011101110111011101110111011101110111011101100110011001100110011001100110011001100101010101010101,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010001000100100001001001000110011001100111011001100111011101100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001100110011001100111011101100111011101100110011001110111011101100110011001100111011101110110011001100110010101010101011001100110011101100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101010101000100001100110100010101010100010001000011001100110011001000100010001000100010001100110011001100110100010001010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100110010001000100010001100110100010001010110010101010101010101010110011001100110011001110110011001110110011001010011001101000011001000100010001000100010001000100010001000110100010000110010001000010001000100010001000100100010001000100010000100100010001000100010001000100010001000100010001000100010001000110100011001110111011101110111011101100110011001010101011001100110011001010101010101010100010001000011001000100010001101000100001101000101010001000100010001000100010001010101011001100101010001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010100110010001000100010001000100010001000100011010000110011010000110010001000010010001000100011001100110011010001000100010001010110011001100110011001110111011101110111011101110111011101110111011101100110011001100110011001100101010101100110011001100101,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110001000100010010001001010110011001100110011001100110011101100111011101100110011001100110011001100110011001100110011001110111011101110111011101110111011101110110011101110111011101110111011101110110011101110110011101110111011101110110011101110110011001100110011001100101011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101100110011001100101010101000100010001000100010001010100010001000100001100110011001100100010001000100010001000110011001101000100010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100100010001100110011001101000101010001100110010101010101011001100110011001100111011101110111011101110110011001100011001100110010001000100010001000100010001000100010001101000101010101000010001000100001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100011001110111011101100111011001100110011001010101011001100110011001100110010101100101010001000011001000100011001101000100010001000100010001000100010001000100010001000101010101010100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010000110010001000100010001000100010001000100011010001000100010001010100001100100001000100100011001101000011010001000100010101010110011001100110011001100111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100101,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001000100010010001101100110011101100110011001100110011001100111011101100111011001100110011001110110011001100111011101100110011101110110011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100101010101010101010101010100010001000101010101000011001100110011001000100010001000100010001000110011001101000100010101010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001000100011001100110100001101010101010101100110010101010101011001100110011101110111011101110111011101110111011101010011001000100010001000100010001000100010001000100011010001000101010100110010000100100010000100010001000100100010001000100011001000100010001000110010001000100010001000100010001000100010001000100011010101110110011101110111011101110111011001010110011001100110011001100110011001100110010101010100001100100011001101000101010101000101010001010101010101010101010101000101010101000011010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010000110010001000100010001000100010001000110011010001010100001101000101010000100001000100100011001101000100010001000100010101010110011001100110011001110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100101,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100001000100010010010001100110011001110110011001100110011001100110011001100110011001110111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010101010101010101010001000100010000110011001100110011001000100010001000100010001000110011010001000100010101010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001100110011001000110011001101000101010001010101010101100110011001100110011001110111011101110111011101110111011101110111011101010011001000100010001000100010001000100010001000100011010001010101010101000010000100010010000100010001000100100011001100110011001100110011001100110010001000100010001000100010001000100010001000010011010101110111011101110111011101110111011001100110011001100110011001100110011001100110010101100101010000110011001101000101010101010101010101000101010101010101010101010101010101000100011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100010000110010001000100010001000100010001000110100010001010101010001000100001100010010000100100011010001000100010001000100010101100110011001100110011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100101,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000010001001000100010010101100110011001110110011001100110011001100110011001100110011001110110011001100110011101100110011001110111011001100110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001010101010101010101010101000100010000110011001100110011001000100010001000100010001000100011001101000101010101000101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000011001100110011001100110011001101010101010001100101011001100110011001100110011101110111011101110111011101110111011101110111011101100011001000100010001000100010001000100010001000100100010101010101010101000010000100010001000100010001001000110011001100110100010001000011001100110011001100100011001000100010001000100010001000100010010101100111011101110111011101110111011101100110011101100110011001100110011001100110011001100110010100110011001101000100010101100101010101010101010101010101010101010101010001000101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100010000100010001000100010001000100011001100110100010101010110010101010101010000100010000100100011010001000100010001010101010101100110011001100110011101100111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100010001000100100011011001100110011001100110011001100111011101110111011101110111011101110110011001100110011001100110011001100110011101110111011101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100101010101010101010101010100001100110011001100110011001000100010001000100010001000110011001101010100010001010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011000110011010000110011001101000100010001010101010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101100011001000100010001000100010001000100010001000110101010101100110010101000010000100010001000100010001001000110100010001000100010101010011010001000100001100110011001100100010001000100010001000100010010101110111011101110111011101110111011101110111011101110111011101100110011001100110011001110110011001010100010000110100010101100110010101010101010101010101010101010101010101000101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010100010000100010001000100010001000110011001100110100010101100110011001010110010000010001000100010010010001010100010001010101010101100110011001100110011001100111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000010001000100100011011001100110011001100110011001100110011001100110011001110110011001110111011001100110011001100110011001100110011001100110011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110010101010101010101010100001100110011001100110010001000100010001000100010001000110011010001000100010001010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000110100010000110011010001000100010101100101010101100110011001110110011101110111011101110111011101110111011101110111011101110111011101100011001000100010001000100010001000100010001101000101011001100110010101000011000100010001000100010001001001000100010101010101010101010100010001000100001100110011001100110011001000100010001000100010010001110111011101110111011101110111011101110111011101110111011101100111011001110110011001110110011001100101010101000100010001100110011001010101010101010101010101010110010101000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000100001100100010001000100011001000110011010001000100010101100110011001100110010000100001000100010010010001010101010001010101011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001001000100100011001100110011001100110011001100110011001110111011101110111011001100111011101110110011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001010101010101000011001100110010001100110011001000100010001000100010001000110100001100110011001100110100010001010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000100010001000100010001000100010101100101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101010010001000100010001000100010001000100011010001010110011001100110011001010011001000010001000100010010001101000101010101010110010101010100010101010101010001000011001100110011001100100010001000100010001101100111011101110111011101110111011101110111011101110111011101100111011001110110011001110111011101100110011001000100010001010110011101100101010101010101010101100110010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000100001100100010001000110011001100110100010001010101011001100110011001100110010000100001000100010010010001010101010001010101011001100110011001110111011101110111011101110111011101110111011101110111011101100111011101110110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100011000100010001001000100101011001100110011001100110011001100110011001110111011001110111011101110110011001100110011001100111011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110010101000011001100110011001100110011001000100010001000100010001000100010001000110011001100110011010001000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101000101010001010100010001000100011001100101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000100010001000110011010101100110011001100111011001010100001000010001000100010011010101010110011001100101011001100101010101010101010001000100010001000011001100100011001000100010001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100010001010110011001100101010101100110011001100110011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100001000100010001000110011001101000100010001010101011001100110011001100110010000100001000100010010010001100101010101010110011001100111011001110110011001110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000100010001001000110110011001100110011001100110011001100110011001110111011001110111011101110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110010100110011001100110011001100100010001000100010001000100010001000100010001000100010001100110011010001000101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010001010100010001010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100100010001000100010001000100010001000100100011001100110011001110111011101100101001000010001000100010011011001100111011101100110011001100110011001010101010101010101010001000100001100110011001000100010000101000111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101100101010001010110011001100101011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001000100010001000110011001100110100010101010110011001100110011001100110010100110001000100010010001101010101010101010110011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010001000100010001001001000110011001100110011001100110011001100110011101110110011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001010100010101000011001100110011001000100011001000100010001000100010001000100010001000100010001100110100010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101010101010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100100010001000100010001000100010001000110110011001100111011101110111011101100101000100010001000100110101011001110111011101110111011101110110011001100110011001100101010101010100001101000011001000100010001000110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010110011001100110011001100110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100011001000100010001000110011001101000101010101010110011001100110011001100110011001000001000100010010001101010110010101010110011001100110011101110111011001110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110001000100010001001001010110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011001100110011001100101010101000011010001000100001100110011001100100010001000100010001000100010001000100011010001010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101100110010101100101010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001000100010001000100010001000100010001101010110011101110111011101110111011101110101000100010001001001000110011101110111011101110111011101110111011001100110011001100110011001010100010001000011001000100010001000100100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010110011001110110011001100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010010001000100010001000110011001101000100010101100110011001100110011001100110011001010001000100010011010001000110010101010110011001100110011101110111011101100111011101110111011101110111011101110111011101110111011101100111011101100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001000100010001001001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010001000100010000110011010001000100010001000011001100100010001000100010001100110010001000110011010001000100010101010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101100101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010001000100010001000100010001000100010001101010111011101110111011101110111011101110100000100010001001101010111011101110111011101110111011101110111011101100110011001100110011001100101010101000011001000100010001000010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000010001000100010001100110011010001000100010101100110011001100110011001100110011001010001000100100010010001000110011001010110011101110110011101100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100010001000100010001101100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010000110011001100110011001100110011001101000011001100110011001000100010001000100010001100100010001101000100010001000100010101010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000100010001000100010010001010111011101110111011101110111011101110011000100010001010101100111011101110111011101110111011101110111011101100111011001110110011001100110010101010011001100100010001000100010001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110010001000100011001100110100010001000101010101100110011001100110011001100110011001100010000100010010010001010110011001100110011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100010010001000100010010001100110011001100110011001100110011001100110011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101000100010001000100010001000100010001000100010001010100010000110011001000100010001000100010001000100010001101000100010001010101010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110110011001100101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100100010001000100010001000100010001000100010010001010111011101111000011101110111011101100010000100010010010001100111011101110111011101110111011101110111011101110111011101110111011101110110010101000011010000100010001000100010001000110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010000100010001000100011001100110100010001000101010101100110011001100110011001100110011001100010000100010010010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101100110011001100110011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000010010001000100011010101110110011001100110011001100110011001100110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101010101010101010101010101010101010101010101010101010100001100110011001000100010001000100010001000100010001000110100010001010100010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010101110111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001000100010001000100010001000100010001000100010010001100110011101110111011101110111011101100010000100010010010001100111011101110111011101110111011101110111011101110111011101110111011101110110010101000101010000100010001000100010001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101001100100010001000100011001100110100010001010101011001100110011001100110011001100110011001100010000100100010010001010110011101110111011101110111011101100111011101110111011101110111011101110111011101110111011001110111011001110111011001100110011001110110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010010001000100011011001100110011001100110011001100110011101100110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101100101010101010101010101010101010101010101010000110010001100110011001000100010001000100010001000100010001000100010001101000101010101010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101100110011001010101010101100111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010001100100010001000100010001000100010001000100010001101100110011101110111011101110111011101010001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110110010001010101001100110011001000100010001000100011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100100001100100011001100110011001100110100010101010101011001100110011001100110011001100110011001100011000100100010010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011001110111011001100110011101100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100011000100010001001000100100011001100110011001100110011001100110011101110111011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010110011001010101010101010100001100110011001100110011001000100010001000100010001000100011001000100010001000110100010101100101011001110111011001110111011101110111011101110111011101110110011101110110011101100110011001100110010101000100010001010110010101000100010001010101010001000101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001100100010001000100010001000100010001000110011001101010110011001110111011101110111011101010001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101100101010101100101001101000011001000100010001000100010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100001100110011001100110011001100110101010101010101011001100110011001100110011001100110011001100011000100010010010001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011001100111011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000100010010001000100101011101100110011001100110011001100110011001100111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110010101000010001100110011001101000011001000100010001000100010001000100011001100110010001100110011001101000110011001100111011001110111011101110111011101110111011101110110011001100111011001100110011001100101010101000100010001000110010101000100010000110011001101000101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000011001000100010001000100010001000100010001000110100001101000110011101110111011101110111011101000001000100010011011101110111011101110111011101110111011101110111011101110111011101110111011001010110011001100100010001000011001100100010001000100010001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100100001100110011001100110011001101000101010101010101011001100110011001100110011001100110011001100011000100010010010001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010010000100010010001000110110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100101001100100011001100110011010001000010001000100010001000100010001000100010001100110011001000110011001100110100010101100110011101100111011101110111011101110111011101110111011001100110011101100110011001100101010001000100010001000101010101000100001100110011001101000100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010100110011001000100010001000100010001000100010001000110100001100110110011101110111011101110111011100110001000100010100011101110111011101110111011101110111011101110111011101110111011101110111010101100111011001010101010001000011001100100010001000100010001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100100001100110011001100110011001101000101011001100110011001100110011001100110011001100110011001100100000100100010010001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101100111011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000001000100100001001001000110011001100110011001100110011001100110011001100111011101110110011101110110011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001000011001100110011001100110011010000110010001000100010001000100010001000100010001000110100001100110011001100110011001101010110011001100111011101110111011101110111011101110111011101100110011001100110011001100101010001000100010001000100010101000011001100110011001101000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010000110011001000100010001000100010001000110011001000110100010001000100011101110111011101110111011100110001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011001110111011001010101010001000100001100100010001000100010001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010011001100110011001100110011001101000101011001100110011001100111011001100110011001100110011001100100000100100010010001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110001000100010001001001000110011001100110011001100110011001100110011001100110011101110110011001110111011001100110011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101100111011101100110011001110110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110010000110011001100110011001100110011010000110010001000100010001000100010001000100010001000110100010000110011001100110011001101000100010101100110011001110111011101110111011101110111011001110110010101010110011001100101010000110100010001000100010000110011001100110011001101000101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100010000110010001000100010001000100010001000110011001100110101010001000100010101110111011101110111011100100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101100101010101010100001100100010001000100010001101000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001000011001100110011001100110011010001000101011001100110011001100111011101110110011001110110011001100011000100100010001101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001000100010010001001010110011001100110011001100110011001100110011001110111011101110110011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101100110011001100110011001100111011101100111011101100111011101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100100001100110011001100110011001100110011001100110011001000100010001000100011001000100010001000110100010000110011001100110011001101000100010001010110011101110110011101110111011101110110011001100111011001010101011001100101010001000011001100110011001100110011001100110011001101000101010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100100010001000100010001000100010001100110011001100110101011001000101010101100111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101010101001100100010001000100010001000110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101000011001100110011001100110011010001010110011001100110011001100110011001100110011101110110011101100011000100010010001101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100001000100100010001101100110011001100110011001100110011001100110011001100110011001100111011101100111011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011001100110011101100110011001100110011101110110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011000110011001100110011010000110011001100110011001100110011001000100010001000110011001000100011001100110100010001000011001100110011010001000100010001010110011101110111011101110111011101110111011001100110011001100101010001010101010001000011001100110011001100100010001000100011001101000101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000011001100100010001000100010001000100010001100110100010000110101011101010100011001100111011101110111011000100001000100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100101011001010101001100100011001000100010001000110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000011001100110011001101000100010001010110011001100110011101110110011101110111011101110110011101110011000100010001001001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000100001000100100010010001100110011001100110011001100110011001100110011001100111011001100110011101100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101100111011101100110011101100110011001100110011001100110011001100110011001100110011001100110011001100101011001100111011001110111011101110111011101110111011101110111011101110111011101110110011001100110010000110011001100110011001100110011001100110011001100100010001000100010001000110011001000100011001100110011010001010100001100110011010001000100010001010101011001110110011101110111011101110111011101100110011001100110010101000100010000110011001100110011001100110010001000110011001101000101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001000100010001000100010001000100010001100110100010001000100011001110101011001110111011101110111010100100001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100001000110011001000100010001000110100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110100001100110011010001000100010001010110011001100110011101110111011101110111011101110110011001110100000100010001001001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100010001001000100011010101100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011001100111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110011001110110011001100110011001100110011001100110011001100110011001100110010101100110011001100101011001100110011001100101010101100110011001100110011101110111011101110111011101110111011101110111011101100110011001010011001100110011001100110011001101000011001100110011001100110011001000100010001000110011001000100011001100110011010001000101010000110011010001000100010001010101011001110111011101110111011001110110011001100110011001100110011001100100001100110011001100110011001100110011001000110011010001000100010101010110011001100110011001110111011101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001100110010001000100010001000100010001100110101010101010101011001110110011001110111011101110111010100100001000101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100001001000011001100100010001000110100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110100010001000100010101010110011001100110011001110111011101110111011101110111011001110100000100010001001001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000010010001000110011010101100110011001100110011001100110011001100110011001100110011101110110011001100111011101100111011101100111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010110011001100110010101010110011001010101010101010110011001010110011001110111011001110111011101100111011101110111011101100110010100110011001100110011001100110100010001000100010000110011001100110011001000100010001001000011001000100011001100110011010001000101010001000100010001000100010001010101011001110111011101110111011101100110011101100110011101100110011001100110010000110011001100110011001000100010001000110011010000110100010001010110011001100110011001100110011001010101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110010001000100010001000100010001101000101011001100110011001110111011001110111011101110111010100010001000101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100011001101000011001100110010001001000100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100001101000100010001010100010101010110011001100110011001110111011101110111011101110111011001110101000100010001001001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000010010001000110100011001100110011001100110011001100110011001100110011001100111011001100110011001100110011001110111011001100111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011001110111011101110111011001110110011001100110011001100110011001100110011001100110011001100110011001100101010101000100010101100110010101000100010101010100010001010101010101000100011001100111011101110111011001100110011101110111011101100101001100110011001100110011001101000100010001000100010001000011001100110011001000100010001000110011001100110011001100110011001101000101010101000100010001000100010001010110011001110110011001100111011101100111011001100110011001100110011001100110010100110011001100110010001000100010001100110011001100110011010001010101010101100101010101100101010101000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110011001100100010001000100010001000100011001101000101011001100110011101110111011101110111011101110111010000010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010011010101010100010000110010001001000101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100001101000100010001010101010101100110011001110111011101100111011101110111011101110111011101110101001000010001001001000110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010010001000110101011001100110011001100110011001100110011001100110011001100110011001110111011101110111011001100111011101110110011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101100111011101110110011001100110011001100110011001100110011001100110011001100110011001010101010001000100010001000101010101010100010001000100010001000101010101000100010101100110011001100110011001100110011101110111011001100100001101000011001100110011010001000100010001010100010001000011010001000011001000100010001000100010001100110011001100110011001101000101010101010100010001000100010101010110011001110111011101110110011001100110011001110111011101100110011001100101001100110011001000100010001000100010001000100011001100110011010001010101010101010101010101010101010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100110010001100100010001100110010001000100011010001000101011001100110011101110111011101110111011101110111010000010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010100011001010100010000100010001101000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000100010001000100010001010101011001100110011001110111011101110111011101110111011101110111011101110110001000010001001001000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100011000100010010001100110101011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110110011001100110011001100110011001100110011001100110011001100110011001010101010001000100010001000100010001010100001100110011010000110100010101000100010101010110010101100110011001100110011001010101011001100101010101000011010001000100010001000101010101010101010101000100010001000011001000100010001000100010001000100011001100110011010001000101010101010101010101000100010101010110011001100111011101110110011101110110011001100110011001100110011001100100001100110010001000100010001000100010001000100010001100110100010101010101010101000100010001010101010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000011001100110011001100110011001100110011001000100011010001000101011101110111011101110111011101110111011101110111001100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101011001010100010000100010001101000101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000100010001000100010001010101011001100110011001110111011101110111011101110111011101110111011101110110001000010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100010000100010010001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101100110011001100110011101110111011101110111011101110111011101100111011101100110011001100110011001100110011001100110011001100110011001100110010101010101010001000100010001000100001100110011001100110011001100110011010001000101010101010101011001100110011001100101010001000101010101100101010000110100010001000100010101010100010101010101010101000101010100110011001000100010001000100011001100110011001100110011010001000101010101100101010101010100010101100110011001110111011101100110011001100101010101000100010001000011001101000100010000110010001000100010001000100010001000100010001100110100010001010100010001000100010101010101010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000101010100110011001100110011001101000011001100110100010001010101011101110111011101110111011101110111011101110111001100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010110011001010101001100100010001000110101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000100010001010100010001010101011001100111011101110111011101110111011101110111011101110111011101110110001100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001010010000100100010001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001110111011001100111011101110111011001100111011001100111011101110111011101110111011001100111011101110111011101100110011001100110011001100110011001100110011001100110011001010101010101010101010001000100010001000100010000110011001100110011001100110011001100110100010001010101011001100110011001000100010001010101011001100101010001000101010001000100010101010101010101010101010101010101010000110011001000100010001100110011001100110011001100110100010001000100010101010101010101100101010101100110011001100111011101100110011001010101010101010100010001000011001100100011001100110011001000100010001000100010001000100011001101000100010001000011010001000100010101010101010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110010000110011001100110011001101000100010001000100010101010110011101110111011101110111011101110111011101110110001100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101100110011001010101001100100010001000110101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000101010001010101010101010101011001100111011101110111011101110111011101110111011101110111011101110111001100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001000001000100100010001101010110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011001110111011001100111011101100110011101100110011101110110011001100110010101100110011101100111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100101010001000100010001000100001101000100010001000011001100110011001100110011001100110011010001010101011001100110010101000100010001010101011001010101010101010101010001010101010101010101010101010101010101010101010000110011001100110010001100110011001100110011001100110100010001000100010101100110010101100101010101100110011001100110011001100110010101010101010101010101010101000011001100110010001000110011001100110010001000100010001000100011001101000011001100110011001101000101010101010101010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010100001100110011010001000100010001010110010101010101011001100110011101110111011101110111011101110111011101110110001000010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010000100010001000110101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001010101010001010101010101010101011001100111011101110111011101110111011101110111011101110111011101110111010000010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011000110001000100100010001101010110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001100110011001100110011001100110011001110110011001110110011101100111011101110111011001110111011101110111011101100110011001100110011001100110011001100110011001100110011001100101010101010100001100110011001100110011010001000100001100110010001100110011001100110100010001010101011001010101010000110100010101010110011001100110010101010100010101010101011001010101010101010101010101010101010000110011001100110011001100110011001100110011001100110100010101000100010101100110011001100110010101100110011101110110011001100110010101010110011001100110010101000011001100110010001000100010001000100010001000100010001000100100001100110011001100110011001101000101010001010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000100010000110011010001000101010001010110011001100110010101100110011101110111011101110111011101110111011101110110001000010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110010101010100010000110010001000110101011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001010110010101010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111010000010001000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110010100100001000100010010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100111011101110111011101100110011001100110011001110110011001110111011101100110011001100110011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000011001100110011001100110100010000110011001000100010001100110011010001010101010101010100010001000101010101100110011001100110010101010101010101010110011001010101011001010101010101010101010000110011001100110011001101000011001100110011010001000100010101010100010101100110011001100110010101100111011101110110011001110110011001100110011001100101010001000011001100110011001000100010001000100010001000100010001000100011001000100011001100110011001101000100010001010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000100010000110011010001010101010101010110011001100110010101100111011101110111011101110111011101110111011101110101001000010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010100010000110010001000110100010101100110011101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111010100010001000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110010100010001000100010010010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001100110011001100110011001100101011001110111011001110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010000110011001100110011001100100011010000110011001000100010001000110011010001010101010001000100010001000101010101100110011001100110010101010101010101010101010101000101010101010101010101010101010000110011001100110011001101000100001100110011010001000100010101010101010101100110011001100110011001100111011101100110011101110111011001100110011001100101010000110011001100110011001000100010001000100010001000100010001000100010001000110011001100110011001100110100010001010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100010000110100010001010110011001010110011001110110011001100111011101110111011101110111011101110111011101110101001000100001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010110010100100010001000100100011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111010100010001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110001100010001000100100011010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110110011001100110011001100110011001100101011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100010001000011001100110011001000100010001100110011001000100010001000110011010001000100010001000100010001000100010101100110011001100110011001100110011001010101010101010101011001010100010101010101010000110011001100110011001101000100010000110100001101000100010101100101010101100111011101100110011001100110011101110111011101110110011001100110011001010101010001000011001100110010001000100010001000100010001000100010001000100011001100100010001100110011001100110011010001010110011001100110011101100111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100010001000100010001000100010001010110011001100110011001110111011001100111011101110111011101110111011101110111011101110101001000100001010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101011001100110010100100010001000100100011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011000100001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110001000010001000100100011011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110110011101110110011001100110011001100110011101100110011101100110011001110111011101110111011101110111011001100110011101100110011001100110011001100110011001100110011001100110011001100110010101000100010001000100010000110011001000100010001000100011001000100010001000110011001101000011001100110100010001000101010101100110011001100110011001100110011001100110010101000101010101000100010101010100010000110011001100110011001101000100010000110011010001000100010001100101010101100110011101100110011001100110011101110111011101110111011101100110011001010100010001000011001100100010001000100010001000100010001000100010001000110011001000100010001100110011001100110011001101000100010101010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010100010001000101010001000100010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110101001000100001010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100110010100100010001000100011011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011000100001000100010100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100101001000010001000100100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110110011001100110011001100110011001010110011001110110011001100111011101100110011001100110011001110110011001100110011001100110011001100110011001100110011001010101010001000101010001000100010001000100001100110010001000100010001000100010001000100010001000100011001100110011001100110100010001010101010101010110011001100110011001100110011001100101010001000100010000110100010000110100010000110011001100110100001101000100010001000100010001000100010001010101010101100111011101110111011101100111011101110111011101110111011101110110011001010101010001000011001100110010001000100010001000110011001000100010001000110011001000100011001100110011001100110011010001000101010101100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010001000101010001000101010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110100001000100010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110010100100010001000100011011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110110011001100110011001100110011001100110011001110110011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010001000011001100110011001100100010001000100010001000100010001000100010001000100011001100110011001101000101010101010101010101010101011001100110011001100110011001010100010000110011001100110100010000110100010000110011001100110100010001000100010001000100010001000100010001010101010101100111011101110111011101110111011101110111011101110111011101110110011001010101010101000011001100110011001000100010001100110011001100100010001000100011001100110011001100110011001100110100010101010101011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010001010101010001010101011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110100001000010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010100110010001000100011011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100011000100010001001000110101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110110011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000100010001000011001100110011001000100010001000100010001000100010001000100010001000100011001000100011001101000101010101010101010101010110011001100110011001100110010001000100010000110011001100110100010001000100001100110011001101000100010001000100010001000100010001000100010001000101010101100111011101110111011101110111011101110111011101110111011101110110011001010101010101000011001100110011001100110011001100110011001100100010001000100011001100110011001100110011010001000101010101010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101100101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110011001000010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111010100110010001000100011010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100010000100010001001000110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100111011001100110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001000100010001000011001100110011001000100010001000100010001000100010001000100010001000100010001000100011010001000100010101010101010101100110011001100110011001100101010000110011001101000100010001000100010001000100001100110011001101000100010001010100010101000100010001000100010001000101010101100111011101110111011101110111011101110111011101110111011101110110011001100101010101010100001100110011001100110011010001000100001100100010001000100010001100110011010001000100010001010101010101010110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101100101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101100011001000010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001000100011010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001010010000100010001001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110010101100110011001100110011001100110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001010100010001000011001100110011001000100010001000100010001000100010001000100010001000100010001100110100010001000100010001000101010101100110011001100110010101010101010001000100010001000100010001000100010001000100001100110011001101000100010001010101010101010100010001000100010001010101010101100111011101110111011101110111011101110111011101110111011101100110011001100110011001010100001100110011001100110100010001010011001000100010001100110011001100110011010001000100010001010101010101010110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101100010001000010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001000110011010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001000010000100010001001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010001000100001100110011001000100010001000100010001000100010001000100010001000100010001100110100010001000100010001010101011001100110011001100110010101010101010001000100001100110011001101000100010001000100001100110011001101000100010001010101010101010100010101000100010001010101010101100111011101110111011101110111011101110111011101110111011101110110011001100110010101000011001100110011001101000100010000110010001000100010010001010100010001000011001101000100010101010101010101010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001010101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001100110011010101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011000110001000100010010001101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101000100001100110011001100110010001000100010001000100010001000100010001000100010001101000100010001000100010001010110011001100110011001100110010101010100001100110100010001000100010001000100010001000100001100110011010001000100010001010101010101010101010101010100010001010101010101100111011101110111011101110111011101110111011101110111011101110111011001010100001100110011001100110011010001000100001100100010001000100010001001000100010101010100010001000100010001000101010101010101010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000011001100110100011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110010100100001000100010010001101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101000011001100110011001000100010001000100010001000100010001000100010001000100011001101000100010000110100010001010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011010001000100010101010101011001100101010101010101010101010110011001100111011101110111011101110111011101110111011101110111011101100101010000110011001100110011001100110100010101000011001000100010001000100010001000100011001100110011001101000100010000110011010001010110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000100001100110100011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110010100100001000100010010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010000110011001100110011001000100010001000100010001000100010001000100010001100100011010001000011001100110011001100110011001100110011001100110011010001010100010001000100010001000100010001000100010001000100001100110011010001000101010101010101011001100110011001010101010101010110011001100111011101110111011101110111011101110111011101110111011001000011001100110011001100110011010001000101010101000010001000100010001000100010001000100010001100100011001100110011010001010100010001000101011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000100001100110100010101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010001000100010001001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110001100010001000100100011010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100010001000100001100110011001000100010001000100010001000100010001000100010001000100010001100110010001100110010001000100011010001010101010001000100010001000100010001000100010001000100010001010100010001000100001100110011010001000101010101010101011001100110011001100110010101010110011001100111011101110111011101110111011101110111011101100101010000110011010000110011001100110100010101010100010000110010001000100010001000100010001000100010001000110011001100110011001101000100010101000011010001010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100001100110100011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110001000010001000100100011010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010001010100001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001010110010101010101010001000100010001000100010001000100010001000100010001000100001100110100010001000101010101010110011001100110011001100101010101100110011001100111011101110111011101110111011101110110010101000011001100110100010000110011001101000101010101000100010000100010001000100010001000100010001000100011001000100011001100110011001101000100010001010100010000110100010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010000110100011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100101001000010001000100100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001000101010101010100001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001101010110011001100110010101000011010001000100010101000100010001000101010001000100010000110100010001000101010101010110011001100110011001100110010101100110011001110111011101110111011101110111011001010100001101000100010001000100001101000100010001010110010101010100001100100010001100100010001000100010001000100010001000110011001000110011001100110011010001000101010101000011010001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010001000101011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100100000100010001000100100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001010110010101010100001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000101011001100110011001010100010001000100010101000100010001000101010001000011010000110100010001000101010101100110011001100110011001100110011001100110011001110111011101110111011101110110010000110011010001000100010001000100010001000100010101010101010101010011001000100010001000100010001000100010001000100011001000110011001100110100001100110011010001010100010101010100001100110100011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010001000101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100011000100010001001000110101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001010100001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010001010101011001100110011001100101010001000100010001000100010001000101010101000011001100110100010001010101010101100110011001100110011001100110011001100110011001100110011101110111011001010100010001000011010001000100010001000100010001000101011001010101011001000011001000110010001000100010001000100010001000100011001100110011001100110100010000110100010001000100010001000100010001000100010001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011000100010001000101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001010010000100010001001000110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010000110010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010101010101011001100110011001100101010101010100010000110100010001000101010101010011001101000100010001010101011001100110011001100110011001100110011001100110011001110111011001110110010001000100010001000100010000110100010001000100010101010110010101010101010100110010001100110010001000100010001000100010001000100011001100110011001100110100010001000100010001000100010001000100010001000100010001000101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001000001000100010001001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100101010100110011001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011010001000101010101100110011001100101010101010100010000110011010001010101010101000011001100110100010001010110011001100110011001100110011001100110011101100110011001110111011001010100010001000100010001000100010001000100010001000101010101010101010101100110010000100011001100110010001000100010001000100010001000100010001100110011001101000011010001000100001101000100010001000101010001010101010101000100010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011000110001000100010001001001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010100010001000100010000110100010001000100010001010101010101000011001000100011001100110011001100100010001000100010001000100010001000100011001100110011001100110011001100110100010001010110011001100110010101010101010000110100010001010101010100110011001100110100010001010110011001100110011001100110011001110110011001100110011001110110010101000100001101000100010001000100010001000100010001010101011001010101010101100101001100100011001100100010001000100010001000100010001000100010001000110011001101000011010001000100010000110100010001000101010101000101010101010101010001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110010100100001000100010010001101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110010101010101010001000011001100110011001100110011001100110011001000100010001000100010001000100011001101000011001000110011010001000100001100110010001000100010001000100010001000100010001000100010001000100010001100100011001100110100010101010110011001100101010101000100010001010101010100110011001100110100010101100110011001100110011001100111011101110111011101100110011001100101010000110011010001000100010001000100010001000101010101010101011001100110011001010011001100110011001000100010001000100010001000100010001000100010001100110011001100110011010001000100010001000100010001000101010101000101010101010101010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110010000010001000100010010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000100001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000100010001000100010001100110011001100100010001000100010001000100010001000100010001000100010001000100010001100110011001000110011010001000101011001100110011001010100010101010101010100110011001100110100010101100110011001100110011001100110011101110111011101100111011001010100010001000100010001000100010001000100010001010110010101010110011001100110011000110011001100110011001000100010001000100010001000100010001000110010001100110011001100110011010001000100010001000100010001000101010101000100010101100110010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101000100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110001100010001000100010010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100101010001000011001100110100010000110011001100110011001100110011001100110011001100110011010000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100100010001000100011001100110011010001000100010001010110011001010100010101010101010100110011001100110100010101100110011001100110011001100111011001100110011001110111011001010100010001000100010001000100010001000100010001010110011001100110011001100101010000110011010000110011001100100010001000100010001000100010001000110011001100110011001100110011010001000100010001000100010001000100010101010100010101010110011001100110010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000010001000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100101001000010001000100010010010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110010101000100001101000100010001000100010001000011010000110011010001000100010101000100001101000101010001000011001100110011001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110100001101000011010001000110011001100101010101010101010100110011001101000100010101100110011101110110011101110111011001100110011101110111010101000100010001000100010001000100010101010100010101100110011001100110011001010100001101000100010000110011001100100010001000100010001000100010001000110011001100110011001100110011010001000100010001000100010001000100010101010100010001010110011001100110011001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000010001000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100100001000010001000100010011010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100101010001000100010001000100010001000100010001000100010001000100010101010101010101010100010001010101010101010100001100110011001100110011001000100010001000100010001100110011001000100010001000100010001000100010001000100010001000100010001100110011010001000100010001000101010101010100010001000101011001100101010101100110010100110011010001000101011001100110011001110110011101110111011101110111011101110110010101000100010001000100010001010101010101100100010101100110011001010100001100110100010001000100010000110011001000110010001000100010001000100010001101000011001100110011001100110011001101000100010001000100010001000100010101010101010001010110011001100110011001100101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100011000100010001000100100011011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001010100010101010100010001010101010101010101010101010101010101010101011001100101010101010100010001010101010101010101010001000100010000110010001000100010001000110011001100110010001000100010001000100010001000100010001000100010001000100011001100100010001000110011001100110100010101010101010101010101011001010100010101010101010000110011010001000101011001100110011101110111011101110111011101110111011101110110010101000101010001000100010101010110011001100101011001110110010001000100010001000100010001000100010000110011001000110010001000100010001000100010010000110011001100110011001100110011001100110100010001000100010001000100010101010101010101010110011001100110011001100101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100010000100010001000100100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001010101010101000101010101010101010101010101010101100110011001100110011001100110011001100100010101100101010101010101010001000100001000100010001000100010001100110011001100110010001000100010001000100010001000100010001000100010001100110011001100100010001000100010001000100011001101000101010001010101011001000011010001010101010000110011010001000110011001100110011001110111011101110111011101110111011101110110010101010101010101010101010101100110011001100110011001100100010001000100010001000100010001000101010000110011001100100010001000110010001000100010010000110011001100110011001100110011001100110100010001010100010001000100010101010101010101010110011001100110011001100101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100010001000100010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110011001100110011001100110011001010010000100010001000100100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100101010101100110010101010101010000110010001000100010001000100011001100110100001100100010001000100010001000100010001000100010001000100010001000110011001100110010001000100010001000100010001000110011001101000101010000110011010101100101001100110100010001010110011001110111011101110111011001100111011101110111011101110110010101010101010101010101011001100110011001100110010101000100010001000011010001000100010001010101010000110011001100110010001000110010001000100010001100110011001100110011001100110011001100110011010001010101010001000101010101010101010101000101011001100110011001100110010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110001100010001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100111011001100110011001100110011001010010000100010001001000110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110010001010101010101010110011001100110011001100110011001100110011001100110011001100110011001100101010101010110010101010101001100100010001000100010001000110011001101000100001000100010001000100010001000100010001000100010001000100010001000100011010001000011001000100010001000100010001000100010001100110011001100110011010001100101001100110100010001010110011001110111011101110111011001110111011101110111011101100110010101100110011001100110011001100111011001110110010001000100001100110011010001000100010101010100001100110011001100100011001100110010001000100010001100110011001100110011001100110011001100110011001101000101010101000100010101010101010101010101011001100110011001010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100010001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100111011001100110011001100110011000110001000100010001001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010110011001100110011001100101010001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110010101000011001100100010001000100011001100110011010001000011001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100100010001000100010001000100010001000100010001000110011010001010100001101000100010001100110011001100110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100101001100110011010001000100010001010101011001100100001101000100001100100011001100110011001000110011001100110011001100110011001100110011001100110011001100110100010101010100010001010101010101010101011001100110011001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010000010001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110011001100110011001100110011000100001000100010010001001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010000110011001000100010001000110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110010001000100010001000100010001000100010001000110011001101010100001100110100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100001100110011001101000100010101010110011001010011001101000100001100100011001100100010001100110011001100110011001100110011001100110011001100110011001100110011010001010101010001010110010101010101011001100110010101010101011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111010000010001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001110110011001100110011001100110010100100001000100010010001101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100001100100010001000100010001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001000100010001000100010001000100011001101000011001100110100010101100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100111011001010100010000110011010001000100010101100110011001000011001101000011001100110011001000100010001000110011001100110011001100110011001100110011001101000100010000110100010001000101010101010110011001010100010101100110010001000101010101010100010001000110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111010100100001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011001110110011001100110010000010001000100010010001101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000011001000100010001000100010001100100011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001100110011001100110100010101100110011001100101010001010110011001100110011001100110011001100110011001100110011001100111011001100111011001000011010001000100010001010101011001110111011000110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001101000100010001000011010001000101010101010101011001010100010101100101001101000100010000110100010001010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010100100001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100111011101110110011001100110001000010001000100010010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010011001100110011001000100010001000100010001000110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000100011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000110011010001000011010001010101011001100111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000011010001000100010101010101011001010101010001100101001101000100001100110100010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011000100001000100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100111011001100110011001100101001000010001000100010010010101100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000110011001100110010001000100011001000100010001000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010101010101010001010110011001100110011001100110011001100110011001100110011001100110011001110111011101100101010001000100001100110011010001010110011001110110010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001010101011001100100010001010100001101000011001101000100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011000110001000100010001001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110110011001100110011001100100000100010001000100010011011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100001100110011001100110010001000100011001000100010001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011010001000100010101100110011001100110011001100110011001100110011001100110011001110111011101110111011101110101010001000011001100110100010101010110011101110110001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011001101000100010001000100010001000011010001010101011001100100001101000011001100110011001101000100010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001110110011101100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110011000110001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101100110011001100010000100010001000100100100011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000011001100110100001100110010001000100010001000100011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110100010001010101011001100110011001100110011001100110011001100110011001110111011101110111011001010100010000110011010001000101010101100111011101110100001100110011001100110011001100110011001100110011001100110011001100110100001100110100010001000011001101000100010001000100010101000100010001000101010101010100001100110011001100110011010001000101010101100111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100110011101110111011101100110011101110110011001100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011000110001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011101100110011101010010000100010001000100100101011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010000110011001100110010001000100011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001100110011001101000100010101100110011001100110011001100110011001100110011001100110011101110110011001000011001100110011001101000101011001100111011101110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000011010001010101010001000100010101000101010001000100010101100100001100110011001100110011010001010101010101100110011001010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011001100110011001100110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001000010000100010010001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001110111011001100110011101000001000100010001000100100101011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100110100010001010100010000110010001100110010001000110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001101000100010001010101010101010101010001010101011001100110011001100110011001100111011001000100001100110011010001000100011001110111011101100011001101000100001100110011001100110011001100110011001100110011010001000100010001000101010101010100010001010110010101010100010001000100010001000100010101100100001100110011001100110100010101010101010101100101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100111011101100110011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100110011101010010000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011001100111011000110001000100010001000100110110011001100110011001100110011101100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001100110100010101010101001100100010001000110011001000110011001100110011001100100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010001000101010101010101010001010101011001100110011001110111011101110111011001000100010000110011010001000101011001110111011101010011010001000100010000110011001101000011001100110011010000110011010001010100010101010101011001100100010001100110011001100101010101000100010001000101010101010100001100110011001101000101010101010101010001010101011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101100111011001100111011101110110011101100110011101110110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011001100110011101010010000100010001000100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100111010100100001000100010001000100110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100001101000100010101010101001100100011001000110011001100110011001100110100001100100010001000100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011010000110100010001010100010001000100010101010110011001100110011001100111011101110111011000110100010000110100010001000110011101110111011101000100010101000100010001000100010000110011001100110011001100110011010001010101010101010110011001100101010001100110011001100110011001010100010001000100010101000011001100110011001101010101010001000100010001000100011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111100010001000100001111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001100111011101110111011101110111011101110110011001110111011001100110011101100110011001110111011101110110011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100010000100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100111010000010001000100010001000101000111011001100111011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001010100010101000100001100110011001100110011001100110100010001000100001100100010001000100010001000100010001000100011001100100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001000100010001010101010101010110011001100110011001100110011001100110010100110100010000110100010101010110011101110111011000110100010101010100010001000100001100110011001100110011001100110011010001000101011001100110011001100101010001010111011001100110010101010101010101000011010001000011001100110011010001010100010001000100010001000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010000111100010000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101110110011101110111011101110111011001100111011101110111011101110110011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100011000100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001110110001100010001000100010001001001010111011001100111011101100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010001000101010101000100001100110011001100110011001100110100010101010100001100100010001000100010001000100010001100110011001100110010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001000100010101000100010001000101010101010110011001100110011101110111011101110111010101000101010101000101010101010111011101110111011000110101010101010101010001000100001100110011001100110011001100110100010101010110011001100110011001100101010001010110011001100110011001010101010101000100010000110011001100110011010001000100010001000100010001010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000011110001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101100110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100011000100010001001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001110101001000010001000100010001001001100111011001100110011001100110011001100111011001100110011001100110011001100110011001100110010101010110011001100110011001100110011001100110011001100110011001100110010101000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010001000101010101010100001100110011001100110011001100110100011001010011001100100011001000100010001000100010001100110100010000110010001001000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010001000100010001000100010001000100010101010101010101100110011101110111011101110111010100110101010101000110011001100111100001110111011000110110011001010101010101000100010000110011001100110011001100110100010101000110011001100110011001010101010001010101010101010101010101100101010101010100010001000011001100110011010001000100010001000100010001000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101100110011001100110011001100111011001100110011101110110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100100000100010001001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001110100000100010001000100010001001101100110011001110111011001110110011001100110011001100110011101110110011101100110011001100110010101010110011001100110011001100110011001100110011001100110011001100110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001000100010001010101011001010100001100110011001100110011001100110100011001010011001100110011001000100010001000100010010001010100010000100010001101010011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000100001100110011001101000100010101010101011001100110011001110111011101110111010101000101011001010110011101110111100001111000010101000110011001010101010101010101010000110011001100110011001100110101011001000101011101110110011001100101010001000101010001000100010001000100010001000011001100110011001100110011001100110100010001010101010101010110011001010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111011101100111011101110111011101110111011101110111011101110111011101110110011101110111011101110110011101110110011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110100000100010001001000010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100011000100010001000100010010010101110111011101110111011101110111011101110110011101110110011101100110011101100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001000100010001000101011001010011001100110011001000110011001101000101011001000011001100110011001100100010001000100010001101010101001100100010001101000100001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011010001000100010101010101011001100110011001110111011101110111010101000110011001010111011101110111100010000111010001000110011001100110011001010101010000110011001100110011001100110101010100110101011101110110010101100101010001000100010001000100010001000100010000110011001100110011001100110011001101000100010101010100010101010110011001100110010101010111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011001110110011101110111011101110111011101110111011101110110011101100110011001100111011101110111011101110111011101100110011101110111011101110111011101110110011001110111011101110111011101110111011101100110011001110101001000010001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001010010000100010001000100010010011001110110011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100010001000100010001000100010101000011001100110011001100110011001101000101011001000011001100110011001000100010001000100010001000110011001000100010001101010101001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010001010101011001100110011001110111011101110111011001000110011001100111011101110111100010000111001101010111011001100110011001100110010001000011001100110011001101000101010100110101011101110110010101000100010001000100010001000100010001000100001100110011001100110011001100110011001100110100010001010101010101010110011001110111011101100110011101110111011101110111011101111000011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111011110000111011101110111011110000111100001111000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011001100111011101110111011101110111011101110111011001110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101100111011001110101001000010001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001000001000100010001000100010011011001110111011101110111011101110111011101110111011101110111011101100110011001100111011001100110011001000110011001100110011001100110011001100110011001100110011001100101010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000101001100110011001100110011001100110100010001000110011001000011001100110011001100100010001000100010001000100010001000100010001101000101010000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001101000100010101010110011001100110011001110111011001010110011101100111100010001000100010000110001101100111011101110111011101100110010101000011001100110011001101000110010001000101011001100111011001010100010001000101010101010101010101000011001100110011001100110011001100110011001100110011001100110100010101010110011001100111011001110110011001110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011110001000011101110111100010000111011101110111100010001000100001111000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101100110011001110111011101110110011101110111011101110111011001100110011001100110001000010001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100111011000110001000100010001000100010101011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001100110011001000110011001100110011001100110011001100110011001100110011001100101010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001010101010001000100001100110011001100110011001101000100010001010110011001010100001100110011001100110011001100100010001000100010010001000010001101000101010000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000100010001100110011001100110011001100110011001101000100010001010110011001110111011001000110011101100111100010001000100010000110010001110111011101110111011101110111010101000011001100110011001101010110010001000101010101010110010101010101010101000101010101010110010100110011001100110011001100110011001100110011001100110011001100110011010001000101011001100110011001110111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011110000111011110001000011101110111011101110111011101110111011101110111011110000111100010001000011101111000011110001000011110000111011101110111011110001000100010001000011110000111011101111000100001110111100010001000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011001110110011001110111011101110111011101110111011101110110011001110111011001100110001100010001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100111010100100001000100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101100110011001010110011001100110011001100110011001100110011001100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010101100101001101000011001100110011001100110011010001000100010101100110011001010100001100110011001100110011001100100010001101000011010100110011010001000100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001000100010001000100011001100110011001100110011001100110011001101000101011001100110011001010110011101110111100010001000100010000101010001110111011101110111011101110110010101000011001100110011001101010110010001000101010101010101010101010101010001000100010001010101001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001010110011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100001110111100010000111011101110111011101111000100001110111100010001000100010001000100010001000011101111000100010001000100001111000011110001000011101111000100010001000100010001000100010001000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101100110011101110111011001110111011101110111011101110111011101110111011101110111011001100110001100010001000100010010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110010000010001000100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101010101011001100110011001100110011001100110011001100110011001100100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001000101011001100100010000110011001100110011001100110011010001010101010101100110011001010100001100110011001101000100010000110010001101010100010100100011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001100110011001100100011001100110100010001000100011001100110011001010110011101111000100010001000100010000100010101110111011101110111011101100110011001000011001100110011010001100110010001000101010101010101011001100101010001000101011001000011001100110011001100100011001100110011001100110011001100110011001100110011001100110100010101000101011001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101010101010101010101010101010011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100001111000011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111011101110111011101110111011101110111011001100111011101110111011001110111011001110110011001110110010000010001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110001100010001000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101010101011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101100110010101000100010000110011001100110011010000110100010001010110011001100111011001010100010001000100010001000100010000110010010001000011001100100011001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100011001100100011001100110011001100110011001100110100010001000100010101100110011001100110011101111000100010001000100001110011011001110111011101110111011101110111011001010100010001000011010101100110001101000101010101010101011001100101010001010110010000110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001010101010001010111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010000100001000100010001001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111,
	2400'b011001100101001000010001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100101011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001000100010000110011001100110011010001000101010101010111011001110111011101100101010101010101010101010101001100100010001100100010001000100010001000110011010001000011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011010001000100010001010100010101100110011001100110011101111000100010001000100001100011011001110111011101110111011101110111011001000100010000110011010101110110001101010110010101100110011001100101010101100100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010101010101010101010101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000011000010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111010100100010000100010001001101100111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011001100110011001100111,
	2400'b011001100100000100010001000100010001001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100101011001100110011001100110011001100110011001100110011001010100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010011001100110011001100110011010001010110011001100111011101110111011101100101010101010110011001010100001000100010001100100010001000100010001000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110100010101000101010101010101010101100110010101100110011001100110011110001000100010001000100001010100011101110111011101110111011101110111011001010100010000110011011010000110001101010110011001100110011101100110011001000011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110100011001100110010101010101010101010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101010101010101010101011101110111011101110111011101110111010101010101010101010101001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111010100100001000100100001001001100111011101110111011101110111011101110111011101110111011001110111011101110110011001110111011001100110011001100110,
	2400'b011001100010000100010001000100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101011001100110011001100110011001100110011001100110011001010100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010001010110010101000100010000110011001100110100010001100110011001100111011101110111011101110110011001100110010101000011001000100010001000100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011010001000101010001000101010001000100010001000100010101100110011001110111011101110111011001100101011001110111011110001000100010001000100001000101011101110111011101110111011101110111011001010101010000110100011110000101001101010110011001110111011101100111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000011001100110100010101100110011001100101010101010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110101010101010101010101110111011101110111011101110111011101110111011101110101010101010101010101010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100010010000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011000100001000100010001001001010111011101110111011101110111011101110111011101110110011001110111011001110111011001100111011001100110011001100110,
	2400'b011101000001000100010001000100010001010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101011001110110011001100110011001100110011001100110011001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010101100110010101000100010001000011001100110100010101100111011101110111011101110111011101110111011001100110010100100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101000011010001010101010101010101010101010101010001000101011101110111011101110111011101110101011001100111011110001000100010001000011100110110011101110111011101110111011101110111011001010101010000110101011110000101001101100111011101110111011101110101010000110011001100110011001100110011010001000011001100110011001100110011001101000100001101000100001101000100010001100111011101110110010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101010101010101010101001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011000100001001000100001001001000111011101110111011101110111011001100111011101100111011101110111011101110111011001100110011001100110011001100110,
	2400'b011000110001000100010001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110110011101100110011001100110011001100110011001000110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000100010001000100001100110100011001100111011101110111011101110111011101110111011001100101001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010001000100010001000100010101000011010001010110011101110111011101110111011101100111011110001000100010001000011000110111011101110111100010001000011110000111011001100101010000110110100010000101010001110111011101110111100001100100010000110011001100110011001100110011010001000011001100110011001100110011001101000100010001000100010001000100010001010111011101110111011001100110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001101010101010101010101010101110111011101111001100110011001100110011001100110010111011101110111011101110101010101010101010100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011000110001000100010001000101000110011101110111011101110110011101110111011101100111011101110111011101100110011001100110011001100110011001100110,
	2400'b011000100001000100010001000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110110011001100110011001100110011001100110011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101000101010101000100010001000100011001100111011101110111011101110111011101110111011001010011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001000011010001000011001100110100011001100111011110000111100001110111011110001000100010001000010101000111100010001000100010001000100010001000011101110101001101000111100010000100010001110111011110001000011101010101001100110011001100110011001100110100010000110011001100110011001100110011001101000101010000110100010001000100010001000110011101110111011101100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011010101010101010101010101011101110111100110011001100110011001100110011001100110011001100101110111011101110111010101010101010101010011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000010001000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011000110001000100100001000100110110011101110111011101110110011101110111011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b010000010001000100010001000100110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001110111011101100111011001100110011001100110010101000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000101010101010100010001010100011001100111011101110111011101110111011101110111010100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001000110011001100110100010001000011001100110011001101000100010001010110011101110111011110001000100010001000100010001000010001011000100010001000100010001000100010001000100001110101010001000111100010000100010101110111100010001000011001100101001100110011010001000011001101000100001100110011001100110011001100110011001100110101011001000100010101010100010001000101011101111000100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010111011101111001100110011001100110011001100110011001100110011001100110010111011101110111011101010101010101010011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000010010000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100100010000100100110011101110110011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110,
	2400'b001000010001000100010001000101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001100111011101110111011101100110011001100111010101000111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100010001100110010101010101010101100101011001110111011101110111011101110111011101110110010101000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001000110011001100110011010001000100010000110011001101000100010001000101011001110111011110001000100010001000100010000111001101111000100010001000100010001000100010001000100001110100001101101000100001110100010110001000100010001000011101100100010000110100010001000011010001000011001100110011001100110100010000110011001100110100011001010100010101010101010101010101010101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101110111011101111001100110011001100110011001100110011001100110011001100110011001011101110111011101110101010101010101001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000010010000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010010000100100101011101110110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100010001001001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110110001101100111011001100111011101110111011001100111010001010111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011101110110010101010101011001100110011001010110011001100110011001100111011101110111011101110111011101110110010100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000110011001100110100010001000100010101010011001101000100010001000101010101100111011110001000100010001000100010000101010001111000100010001000100010001000100010001000100001110100010001111000100001110100011010001000100010001000100001100101010000110101010001000100010000110011001100110011001100110100010001000100001100110011010101010101010101010110010101010101011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101011101110111011110011001100110011001100110011001100110011001100110011001100110011001100101110111011101110101010101010101010100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000010010000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101010010000100010001000100100100011101110110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100010010001101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001101010111011001100111011101110110011001110110010001010111011101110110011001100110011001100110011001100110011001100110011101110110011001110111011101100101010101010110011001110111011001010110011001110111011101100111011101110111011101110111011101100101001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010001000100010101100100001101000100010001000100010101010110011001111000100010001000100010000100010110001000100010001000100010001000100010001000100001100011010110001000100001100100011110001000100010001000100001100101010101010110010001000100010000110011001100110011001101000100010001000100001100110011010001100110011001110111011101100110011101010110100010001000100010001001100010001000100110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111010101010101010100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111010100100010000100100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101010010000100100010001000100100011101110110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110,
	2400'b000100010001000100100010010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011001100110010001010111011101110111011101100110011001110110010001100111011101110111011101110111011101100110011001100110011001100110011001100111011101110111011101110110010101100111011101110111011001100110011001110111011101110111011101110111011101110111011001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001010100010101010101010101000100010101010101010101010101010101100111100010001000100001110011011010001000100010001000100010001000100010001000100001010011011110001000100001010100011110001000100010001000100001110110010101100110010101010100001100110011001100110011001101010101010001000100010000110011001101010110010101111000011101110110011101100110011110001000100010011000100010001000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010111011101110111100110011001100110011001100110011001101110111011101110111011101110011001100110011001011101110111010101010101010101010011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100110010100100010000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001100110011001100110011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100010000100100010001000010011011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100100010011001100111011101110111011101110110011101110111011101110111011101100110011101110111011101110111011101110110011001110111011101110110010001000111011101110111011001100110011001110101010001100111011101110111011101100111011101110110011001110111011101100111011101110111011101110111011101110110011001110111011101110111011001100111011001110111011101110111011101110111011101110110010000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000100010101010100010101010100010101010110011001100101010101010110011001111000100001010011011110001000100010001000100010001000100010001000100001000100100010001000100001010100100010001000100010001000100010000111010101110110011001010011001100110011010001000100010001010101010101010100010000110011001101010111011001101000011110000111011101110101011010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101110111011101111001100110011001100110011001100110011011101110111011101110111011101110011001100110011001011101110111011101010101010101010011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100110011101100111010100100010000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100011000100010010001000010011011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100100100011001100111011101100110011001100111011101100111011101100111011101100111011001100111011101110111011101100110011001100101010101010110010001010111011101110111011101110111011001110101010001110110011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110101001100110011001000100010001000100010001000100010001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001010101011001100101011001100110011101110110011001100110011001101000100001000100011110001000100010001000100010001000100010001000011101000101100010001000100001000101100010001000100010001000100010000111010101110111011101100011001100110100010001000100010001100101010101010101010001000100001101000111011101101000100010001000011101110101010101101000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101110111011101111001100110011001100110011001100110111011101110111011101111011011100110111011101110011001100101110111011101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011001110111011001110111011101110111010100100010000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110110011001110111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011001000010010001000100010011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100100101011001100110011101100111011101110111011101110111011101110110011001100110010000110100010101100111011001100110011001000011001100100100010101010111011001110111011101100110011001110100010101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101010100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110101011001100101011001110110011101110111011101110110011001100110011000110110011110001000100010001000100010001000100010001000011000110111100010001000100001000110100010001000100010001000100010000111011001100111011101000100010001000100010001000101010001100101010101010101010101000100001101000111100001111000100010001000100010000110010101011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101110111011101111001100110011001100110011001100110011011101110111011101110111011101111011101110111011001100101110111011101110101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011001110111011001110111011101110111011101110111010100100010001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000010010001000100010010101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110,
	2400'b000100010001000100100100010000110110011001100110010101110111011001110111011101110111011001100101001100110011001100110100010101100110011000110011001100110011001101000110011101110111011101100110011101100100011001110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101100101001100110010001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001010110010101110111011101110111011101110111011001100110010100110111011101111000100010001000100010001000100010001000010101000111100010001000100001000111100010001000100010001000100010000111011001010101010101000101010001000101010101000101010101100101010101100101010101000100010001000110100010001000100010001000100110000111010101011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001101010101010101010101011101110111011101111001100110011001100110011001100110111011110111011101110111011011101111011101111111111011100101110111011101110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100110011001110111011101110111011101110111011101110111011101100110010100100010001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001100101001000010001001000100010010101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b000100010001000100100010001100110100001101000011001101010111011001100101010101010110011001100011001000110011001000100010001001000101011001010010001000110011001000110101011001010101010101100110010101000011010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100001100110010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110101011001110111011101110111011101110111011101110111001101000111011101110111100010001000100010001000100010001000010001011000100010001001011101000111100010001000100010001000100010001000011101100101010001010110010001000101010001010110010001010101010101100101010101010100001100110110100110001000100010001000100110010111010101011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001101010101010101010101011101110111011101110111100110011001100110011001100110111101101110111011110111011011101110111101111111011011100101110111011101110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110011001110111011101110111011101110111011101110111011101110111011101100111010100100010000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110001100010001001000100010010001110110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011101110110,
	2400'b000100010001000100100010001000100010001000100011001100110110011001010010001100110011010101010011001000100010001000100010001000100010001101000010001000100011001000100011001100110011001101000100001100100010010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000100001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000100001100110011010001010111011101110111011101110111011101110111001101010111011101110111011101110111100010001000100010000111001101101000100010001001011001001000100010001000100010001000100010001000011101100101010101010110010001000100010101110111010001010110011001010110011001010100010000110110100110001000100010001000100110010111011001011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101011101110111011101110111100110011001100110011001100110111101110110111011110111111101101110011011101110111001100101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101100111010100100010000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100010010001000100010010001100110011001100110011001100110011001100110011001100110011001100111011001100110011101110110011101100110,
	2400'b000100010001001000100010001000100010001000100010001100110011010001000010001000100010010000110010001000100010001000100010001000100010001000110011001000110010001000100010001000110010001000110011001100110011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000011001100110011001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100010001000100010001000101011101110111011101111000100010000110001101100111011101110111011101110111011101111000100010000110001101111000100010001001010101011000100010001000100010011000100010001000100001110110011001100110010001000100011110001000010001111000011101100111011001100101010001000110100110001000100110001001100110011000011101101000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101011101110111011101110111100110011001100110011001100110011011101110111001100111011101101110011001100110011001100101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101100111010100100010000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100100010001000100010001101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111,
	2400'b000100010001001000100010001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100011001100100100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000011010000110010001000100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001101000100010001000100010001000100010001000100010101111000100001110111100010000101001101110111011101110111011101110111011101110111100010000101010001111000100010001000010101101000100010001001100110011001100010001000100001110110011101110110010001000110100010000111010101111000100010000111011101100101010001000101100110011001100110011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110011001100110111011100110011001100110011001100101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100100010001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000100001001000100010001101100111011001110111011001100110011001100110011001100110011001100110011001100110011001110111011001100110,
	2400'b000100010001001000100010001000100010001000100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000110101011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100001100110010001000100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100011001100110010001101000100010001000100010101000100010001000100010001101000100010001000100001110011010101110111011101110111011101110111011101110111011101110100010101110111011110000111010001101000100010001000100010011001100010001001100010000111100010000110010001001000100010000111010110001000100010000111011101110101010101000110100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100010001000100010001000100010001000100010001000100010000111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100100001001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100001000100100010001001010111011001100110011001110110011001100110011001100110011001100110011001100110011101110111011001110111,
	2400'b000100010001001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000110100011001100101010001010100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001101000101010101010101010101010100010001000100010001010111100010001000100001110011011010001000100010001000011110001000011101110111011101100011010101110111011101110110010001111000100010001000100010001000100010001000100010001000100010000110001101101000100010000110011010001000100010001000011101110110010101010110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001100010001000100010001000100010001000100001110111011101110110011001100110011001100111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100100010001000010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010100100001001000100010001001010111011001100110011001100110011101100110011001100110011001100111011001100110011101110111011001110111,
	2400'b000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010101000100010001000011001000110011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101000100001100110011001100100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110100010101100110011001010101010101010100010001010101011110001000100001010011011110001000100010001000100010001000011101110111011101010011011001110111011101110101010001111000100010001000100010001000100010001000100010001000100010000101010001111000100010000101011110001000100010001000100010000111011001100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001011101111001011101110111011101110111010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000011101110111011001100110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000110001000100100010001001000110011001100110011001110110011101100110011001100110011001100110011001110111011101110111011101110111,
	2400'b000100010010001000100010001000100010001000100010001000100010001000110010001000100010001000110011001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100101010001000101010000110011001000100100010101010110010101000100010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101000011001100110100001100110011001000100010001000100010001100100010001000100010001000100010001000110010001000100010001000110011010000110010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011010001100110011101100110011001100101010101010101011010001000100001000100100010001000100010001000100010001000100010001000100001010011011101110111011101110101010001111000100010001000100010001000100010001000100010001000100010000100010110001000100001110101100010001000100010001000100010000111011101110110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011010101010011001101010101001100110011001100110011010101010101010101010101010101010101011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000100100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011001110111011001100111011101110110011001100110011101100110011001100110011001100110011001100110011001100110011000110010000100100010001000110110011001100110011101100111011101110110011001100111011001100110011101110111011101110111011101110110,
	2400'b000100010010001000100010001000100010001000100010001000100010001000100011001100100010001000110011001000100010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001000100010001000100011001000110011001100100010001100110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101000011010001000100001100110011001000100010001000100011001100110010001000100010001000100010001100110010001000100010001101000100001100100010001000110010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001101000110011101110110011101110110011001010101010101111000011100110101100010001000100010001000100010001000100010001000100001000100011101110111011101110100010110000111100010001000100010001000100010001000100010001000100001110100011110001000100101100101100010011001100010001000100010001000100001110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101111001100110011001100110011001100110011001100110011001100101110111011101110111011101110111011101110111010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010000111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001110110011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000100100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001110111011101100110011001100110011001100110011001100110011001000010001000100010001000110110011001100110011001100110011001100111011101110111011001100111011101110111011101110111011101110111,
	2400'b000100010010001000100010001000100001001000100010001000100010001000100011001100100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010100010101010101010000110010001000100010001000110011001100110010001000100010001000100011001100110010001000100011010001000011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011010001000100010000110011001100110101011101110111011101110111011001010111011001011000010100110110100010001000100010001000100010001000100010001000011100110101100001110111011101110011010110001000100010001000100010001000100010001000100010001000100001100100100010011000100001010111100110001001100110011001100110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101111001100110011001100110011001011110011001011101110111011101110111011101110111011101110101010101010101010101010011001100110011001100110011001100110011001100110011001100010000111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110110011001100111011101100111011001100110011101100111011001100110011001100110011001100110011101010010000100100010001000100101011101100110011001110110011001100111011101100111011101110111011101110111011101110111011101110111,
	2400'b000100010010001000100010001000100010001000010010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101000101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101011001100110010000100010001000100010001000110100010000110010001000100010001000110100010000110010001000100100010101000011001000110010001000100010001000100010001100110010001000100010001000100010001000100010001100110011001100110011010000110100010001000100001100110011010101100111011101110111011101100110011001100111010000110111100010001000100010001000100010001000100010001000011000110110100010001000100001110011011010001000100010001000100010001000100010001001100010001000100001000110100010001000011101001000100110001001100110011001100110011000100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101111001100110011001011110010111011101110111011101110111011101110111011101110111011101110111010101010101010101010011001100110011001100110011001100110001000011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001001000010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110110011101110111011101110111011001100110011001100110011001100011000100100010001000100101011001100110011001110111011101100111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100100010001000100010001000010010001000100010001000100010001000110010001000100010001000100010001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101000100010101000100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110110001100100010001000100010001000110011001100110010001000100010001101000100001100100010001001000101010000110011001100110010001000100010001000100010001100100010001000100011001000100010001000100010001000110010001100110100010001000011010001000100001100110011001101000110011101110111011101110101011001010100001000110111100010001000100010001000100010001000100010001000010100110111100010001000100001100011011110001000100010001000100010001000100010001000100010001001011101000111100010001000011001011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101111001100110011001011101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110011001100110011001100010000111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110110011101110111011101110111011001110111011101110110011001110111011001100110011001100011001000100010001000100100011001100110011001100111011101110110011101110110011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100100001100100010001000100010001000110011001000100010001000100011001101010100001100100010001101000100001100110011001100110010001000100010001000100010001100100010001000100011001000100010001000100010001000100011001100110011010001000100010001000100010000110011010001000101010101100111011110000111010101010011001001001000100010001000100010001000100010001000100010001000010001000111100010001000100001010100100010001000100010001000100010001000100010001000100010001001011001001000100010001000010101101001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110011000100001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001001000010011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011001100100001000100010001000100011011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100100001000100010001000100010010001000100010001000100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011001100110011001100100010001100110011001100110010001000100100010101010100001100100011010001000011001101000011001100100010001100100010001000100010001100110010001000100011001100100010001000100010001100110011001100110011001101000100010001000100010001000100010000110100010001000101011001110111010101010011001101011000100010001000100010001000100010001000100010001000001101011000100010001000100001000101100010001000100010001000100010001000100010001000100010011000010101011000100010010111010001111001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010011001100001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010011011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110101001000010010001000100010011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000010001000100010010001000100010001000100010001000010001001000100001001000100010001000100010001000100010001000100010001000100010001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001100100011001100110011001100110010001100110101010101010100001100110011010000110100010001000100001100110011001100100010001000100011001100110010001000100011001100100010001000100010001100110011001100110011001100110100010001000100010001000100010001000100001101000100010001100101011001000011001101111000100010001000100010001000100010001000100010000111001101101000100010001000011101000110100010001000100010001000100010001000100010001000100010000111010001101000100010000110010110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101001100001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110101001000010010001000100010010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000011001100110011001100100011001101000100001100100010001101000110011001010011001100110100010001000100010001000100010000110011001100100010001000100011001100110010001000110011001100100010001000100010001100110011001100110011001100110100010001010101010001000100010101000101010001000100010001000100011001000010001101111000100010001000100010001000100010001000100010000110001101111000100010001000011100110110100010001000100010001000100010001000100010001000100010000110010001111000100010000100011010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010100110000111011101110110011001100110011001100110011001100110011101100110011001100110011001100110011001100110011001100110011001100110011001100111011101110110011001100110011101100111011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010010011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000100001001000110011010001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100100010001000100010001000100010001000100010001000100010001000010001000100010010000100010010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010001000100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000011001100110100001100110011010101010100001100110010001101100110011001000011001101000100010001000100010001000100010000110011001100100010001000110011001100110010001000110011001000100010001000100010001000110011001100110100001100110011010001010101011001010101011001010101010101000100010001000100010000110011010010001000100010001000100010001000100010001000100010000101010001111000100010001000011000110111100010001000100010001000100010001000011101110111011101110100010101110111100001110100011110001000100010001000100110011001100110011001100110011001100110011001100110011001100010001000011101111000100010001000100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101001100110001000011101110111011101110111011101110110011101100110011001100110011101110110011001110111011101100110011101100110011101110111011001100110011101110111011101100111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001001000100010010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100010010001000100010001101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001001000100010001000010001000100010010001000100010001000100010001000100010001000100010000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001100110011001101000100010001000011010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101000011001100110100001100110011011001100101001100110011010001100110010100110011001101000101010101010100010001010100010001000100001100100010001000110011001100110010001000110011001000100011001000100010001000110011001100110100010000110011010001000101010101010101011001100101011001010101010001000100010100110011011010001000100010001000100010001000100010001000100010000100010110001000100010001000010101001000100010001000100010000111011001100110011001010101010101010100010101100110011001010101011101111000100010001000100110011001100110011001100110011001100110011001100110000111011101111000100001111000100010001000100010001000100110011001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110101010100110011000100010000111011101110111011101110111011101110111011101110111011001100110011001100110011001100111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010010010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000010001001000010010001101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000010001000100010001001000100010001000100010001000100010001000100010001000110011001100110100010000110011001101000110011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010100010001000101010000110011011001100101001100110011011001110110010100110011010001010101010101010101010101010101010101010100001100100010001000110100001100110010001000110011001100100011001000100010001000110011010000110100010001000100001101000101010101010110011001100110011001100110010101000100010100110011011110001000100010001000100010001000100010001000100001110011011010001000100010001000010001001000100010001000100001110110011001010110010101010101010101010100010101010101010101000101011001100111011101111000100010011001100110011001100110011001100110011000100001110111011101110111011110001000100010001000100010001000100010011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111010100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010010010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000010001000100100010001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010000100010010000100010010001000010010001000100010001000100010001000100010001000010010001000100010001000100010001000100001001000100010001000100010001000100010001000100010000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110101010101010110010000110100011001100100001100110101011101100110010000110011010001010101010101010101010101010101010101010100001100110010001100110100010000110010001000110011001100100010001000100011001000110011001100110100010101000101010001000100010101010101011001100111011001100111011001010101010000100100100010001000100010001000100010001000100010001000100001110011011010001000100010000111001101011000100010000111011001100110011001100110010101010101010101010100010101010101010101010101010101010101011001100111011101111000100010001001100110011001100010000111011101110111011101111000011101111000100010000111011110001000100010001001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111010100110001000100010001000011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100100001000100010010001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010010001000100010001000100010001000100010001000100010000100010001001000100001000100100010001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100011001100110011001100110011010001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111001100110100011101010011001101000110011101100101001100110100010101010101010101010101011001100110011001010101010000110011001101000101011001000010001100110011001100110011001000100011001100110011010001000100010001010101010101010101010101010110011001100111011001010110011101110110001100110110100010001000100010001000100010001000100010001000100001100011011110000111100010000101001101100111011101100110010101010101010101010101011001010101010101000100010101010101010101010101011001100110011001100101011001100110011001110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111100010001000100110011001101010101001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110101010100110011000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010000100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100100010001001000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010010000100010001000100100010001000100010001000100010001000100010001000100010000100010001001000100010001000010001001000100010001000100010000100010010001000100010001000010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100011001101000101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000110100011001000011001101100111011101100100001100110100010101010101010101010101011001100110010101010100001100110010010001100111011001000010001100110011010000110011001100100011001100110100010101010101010001010101010101100110011101110111011110000111011101010101011101110101001100110111100010001000100010001000100010001000100010001000100001010100011101110110011001100100001101010101010101010101010101010101010101010101010101010101010101000101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111100010001000100010001001100110001000011110000111011110001000100110011001100110011001100110011001100010001001101010101010101010101010101010101010101010101010101010101010101010101011101010111011101110111001100110001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010001001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100001000100010010001000110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100100010000100010010001000100010001000100010001000100010001000100010001000100010000100100010000100010001001000100001000100100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010010001000100010000100010010001000100010001000100010001000110011001101000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000100011010000110011010001110111011001010011001101000101010101010101011001010101010101010101010101010100001100110011010001100110011001000010010001010100010000110011001100110011001000100100011001100110011001100111011001111000100010001000100010001000011101100101011101110100001101000111100010001000100010001000100010001000100010001000100001000100010101010101010101010011010001010101010101010101010101010101010101100101010101010101010101000101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001111000100010011010101010101010101010101010100110101010101010101010101010101010101010101010101010000111011110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110001000100010001001000110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100100010001000100010001000100010001000100001000100100010000100010010001000100010001000100010001000010001001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001100110011001100110100011101110111011101110111011101110111011101110111011001100101011101110111011101110111011101110111011101111000011101110110001100100010001100110011011001110111011001000011001101000110011001100101010101010101010101000101010101000100001100110011010001010110011101000010010001010101010000110011001100110011001100110100011001110111011101110111100010001000100010001000100010001000100001110101010101100011001101011000100010001000100010001000100010001000100010001000011100110100010101010101010101000011010101010101010101010101010101010101011001100101010101010101010001000101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100110011001100010001000100010001000100110011000100110011001100110011001100001110111100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010010001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010000100010001001000100010000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001101000111011101110111011101110111011101100110011001010101010000110100011001110111011101110111011101110111011101110111011101110110001100100011001100110100100001100110010000110011001101010111011101100110010101010101010101010101010101010100001100100011010101100110011101000010010101010100001100110011001100110011001100110100011101110111011110001000100010001000100010001000100010001000100001110110010101010011001101101000100010001000100010001000100010001000100010001000010100110101010101010101010101000011010101010101010101010101010101010101010101010101010101010101010001010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010010001000100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000010001000100010010000100100010000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100011010001100111011101100110010101010100010001000011001100110011001000100011010001100111011101110111011101110111011101110111011101110101001100110011001100110110011101010101001100110011010001100111100001110110010101010101010101100110010101000100001100110011010001100110011001000010010001010100001100110011001100100011001100110100011101110111011110001000100010001000100010001000100010000111011101100110010101000011010001111000100010001000100010001000100010001000100010001000010000110101010101010101010100110100010101010101010101010101010101010110010101010101010101100101010001010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011110001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010000100010010001000100100011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000010001000100010001001000100001000100010010001000100010000100010010001000100010001000100010000100100010001000100010001000010010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100011010001010100010000110011001000110010001100100010001000100010001000100010010001100111011101110111011101110111011101110111011101110101001100110011001101010110010101010100001100110011010101100110011001100101010101010101011001100101010101000100001100110011010001010110011000110010010101010011001100110011001100110011001100110100011001100110011110001000100010001000100010000111011101110111011001000101010100110011010110001000100010001000100010001000100010001000100010000111001101000110010101010101010100110100010101010101010101010101010101010110011001010101010101010101010001010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001110111011101100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010001000100010001000100011011001110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100001001000100010000100100010001000100010001000100010001000100010001000100010000100100010001000100001000100010001001000100010001000100010001000100010001000010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000110011001100100010001000100010001000100010001000100010001000100010000100100011001101000110011101110111011101110111011101110111011101110100001100110011010101010101010001000011001100100100010101010101010101010101010101000100010101010100010101000011001100110011010001010110010100110010010001000100001100110011001100110011001100110100010101010101010101100111011101110111011101110110010101010101010101000101010100100011011010001000100010001000100010001000100010001000100001110101001101010110010101010101010000110101010101010101010101010101010101100110011001100101010101100101010001010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001001001000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011001000100010001000100011011001110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010000100010001001000100010001000100010001000100001000100010010001000100001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100001000100010001000100010001000100100010000100010001000100010001001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001010110011101110111011101110111011101100011001000110100011001010101010000110011001000110100010101010101010101010101010101010100010101000100010101000011001100110100010001010101010000100010010001000011001100110011001100110011001100110011010001010101010101010101010101010101010101010110010101010101010101010101010000100011011010001000100010001000100010001000100010001000011101110101001101010101011001010101001100110101010101010101010101010101011001100110011001010101011001100100010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111100001110111100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001000010001001000100010010101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010000100100010001000100001000100010001001000010001000100010010000100010001001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001010110011101110111011101010011001000100100010101010100010000110011001000110101010101010101010101010101010101010100010001000100010001000011001100110100010001010101010000100010010000110011001100110011001100110011010001000011010001010101010101010101010101010101010101010101010101010101010101000100001100100100011001100111011101111000100010001000100001110111100010000101001101100101010101010100001101000101010101010101010101010101011001100110011001100110011001010100010101100101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111100010001000011110001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001000010001000100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001000010001001000100010010101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100001001000010001000100010001001000100001000100100001000100010001000100100010001000100010000100010010001000100010001000100001000100100001000100010010001000100001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011010101100110011001010011001000110100010101010100001100100010001101000101010101010101010101010101010101010101010101010101010001000011001100110100010101010101010000100011010001000100001100110011001100110011010001000011010001010100010001010101010101010101010101010101010101010101010001000100001100110100010001010110010101010111100010000111011001100111100010000100010001010100010001000100001001000101010101010101010101100101011001100110011001100110011001010100010101100101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000010001000100110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000010001001000100010010001100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001001000100010001000010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010000100010001000100100010000100010001000100100010001000010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101010101010101000010001000110100010101000100001100110010001101010101010101010101010101010101010101010101010101010101010101000011001100110100010001000101010000100011010001000100010000110011001100110011010001000100010001010100010001010101010101010101010001010101010101010100001101000011001100110100010001010101010101000101011101110110010101010101011001100011010001010100010001000011001101010101010101010101011001100110010101010110011001100110011001010101011001100110010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000100010001000110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000100001001000100010001101100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001001000100010000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100010010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001100110100010100110010001000100100010001000011001100110011001101000101010101010101011001010101010101010101010101010101010101000011001101000100010101010101010000100011010001000101010000110011001100110011010001000100010001010101010101010101010101010101010001000100010001000100001100110011001100110100010001010101010001000101011001010100010001000100010001000011010001000100010001000011001101010101010101010101010101010101010101010101011001100110011001000101011001010110010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011110001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000100010001000110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100010010001000100010001001100111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010010001000100010001000100010001000100010001000010001000100010001000100010001000100010010001000100001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001101000100010000110010001000110101010101000010001100110011001101010101010101010101010101010101010101010101010101010101010101000011001101000101010001000100010000100100010101010101010101000100001100110100010101010100010001010101010101010101010101010100010001000100010001000100010000110011001100110100010001000100010001000100010101000100010001000100010000110011001100110100010000110010010001010101010101010110010101010101011001010100010101100110010101000101010101010101010001010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011110001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000010010001000100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100100010001000100010001001010111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010010001000100010001000100010000100010001000100010001000100010001000100010010001000100001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100001100100010001001000101010100110011001100110011010001010101010101010101010101010101010101010101010101010101010101000011001101000101010001000100001100100100010101010101010101000100010001000100010101010101010001000101010101010101010101000100010001000100010001000100010000110011001101000100010001000100010001000100010001000100010001000100010000110011001100110011010000110011010001000100010101010101010101010101011001010100010001010101010001000101010101000100010001000101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101110111011101110111011110001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000010010000100100101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000100010001000100010001001010111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000110100010000110011001100110011010001010101010101010101010101010101010101010101010101010101010000110011010001010100010001000101001100100100010101010101010101010101010001000100010001010101010001000100010001000100010001000100010001000100010001000011001100110011001101000100010001000100010001000100010001000100010001000100010000110011001100110011001100110011010001000100010001000100010001010101010101010100010101010101001101000101010101000100010001000101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101111000011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000010001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100100010001000100010000101000111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000010010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100100001000100100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001001000010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100001100110011001100110011010001010101010001010101010101010101010101010101010101010101010100110011010001010100010001010100001100110101010101010101010101010101010101000101010101010100010001000100010000110011001101000100010001000100010000110011001100110011001101000100010001000100010001000100010001000100010001000100010000110011001100110011001100110011010001000100010001000100010001010100010101010101010101010100010001010101010100110011001100110100010001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100010001000100010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000100010000100110110011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000010001000100100010001000100010000100010001000100010001000100010001000100010001000100010001000100010010000100010001000100010001000100010001000100010001000100100010001000100010001000010001001000010001001000100010001000100010001000100010000100010001000100010001001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100001100110011001100110011010001000100010101010101010101010101010101010101010101010101010000110011010001000011010001000100001100110101010101010101010101010101010101010101010101010100010001000100010000110011001100110100010001000100010000110011001100110011001100110100010001000100010001000100010001000100010001000100001100110011001100110011001100110011010001000100010001000100010001000100010001010100010001000011010001010100001100110011001100110011010001000101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101111000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111001100010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000100010001000100010000100100110011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010010001000010010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100010010000100100001000100010001001000100010001000100010000100010001000100010001001000100010001000100010001000010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100100011010001000101010101010101010101010101010101010101010101010101001100110011001100110011001100110100001000110101010101010101010101010101010101010100010001000100010001000100010000110011001101000100010001000011001100110011001100110011001100110100001101000100010001000100010001000100010001000100001100110011001100110011001100110011010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011010001000100010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110000111011101110111011101110111011101110111011101110111011101110111011101110111001100010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110010001000100010000100100101011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010000100010001001000100010000100010001000100010001000100010001001000100010001000100010001000010001000100010001000100100001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000110011010000110011001100100011010001000100010001010101010101010101010101010101010101000100001100110011010001000100001100110011001000110100010101010101010101010101010101000100010001000011001100110100001100110011001101000011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000011001100110011001100110011001100110100010001000100010101010100010001000101010001000011001100110011001100110011001100110011001100110011001100110100010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011001110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100001110111011101110111011101110111011101110111011101110111011101110111001100010001000100010100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000100010000111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010001000100010000100010100011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100010010001000100001000100010001000100010001000100010001000100010010001000100010001000100010001000100001000100010001001000100010000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001101000011001000100010001101000100010000110011001100110011010001000100010001000100010001000100001101000100010001000011001000110100010001000100010001000011001000110100010001000100010101010101010101000100001100110011001100110011001100110011001101000100010001000011001100110011001100110011001100110100010000110011001101000100010001000100010001000011001100110011001100110011001100110100010001000100010001010100010001000100010001000011001100110011001100110011001100110011001100110011010001000100010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100101010001000100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100110011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000011110001000011110000111011101110111011101110111011101110111010000010001000100010011011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011110000111011101110111100010000111011101111000011101111000100001110111011101110111011101110111011101110111011101110111011101110111011110000111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000010001000100010000100010011011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010010001000100001000100010001001000010001000100010001000100010001000100010001000100010010001000100010001000100010001000010001000100010010001000100010000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100011001101000010001000100010010001000011001100110011001100110100010001000100010001000011001100110011001101000101010101000011001101000100010001000011001101000011001000110100010001000100010001010101010001000100001100110011001100110011001100110011001101000100010001000011001100110011001100110011001100110011001100110011010001000100010001000100001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000011001100110011001100110011001100110011001100110011010001010101010101010101010101100110011001100110011001100110011001100110011001100110011001010110011001100110010101010110011001010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110010101010110011001100110011001100110011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111010000010001000100010011011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100001110111100010001000100010001000011101111000100010001000011110001000011101110111011101110111011101110111011110000111011101110111011101110111100001111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010001000100010001000010011011001110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000010001000100010001001000010010000100010001000100010001001000010001001000100010001000100010001000100010001000100010001000100010000100100010000100010010000100010010001000100001000100010001001000100010001000100010001000100010001000100010001000100010001000100011010000110010001000100010010001000011001100110011001100110100010001000011001100110100001100110100010101010101010000110010001101000100010001000011001101000011001001000100010001000100010001000100010001000100001100110011001100110011001100110011001101000100001100110011001100110011001100110011001100110011001100110011001101000100010000110011001100110011001100110011001100110011001100110011010000110011010001000100010001000100001100110011001100110011001100110011001100110011001100110100010001000100010001000101010101100110011001100110011001100110011001100110011001100110011001010110011001100110011001010110011001100101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001010101011001010101010101100110011001100101010101010101011001110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011110000111011101110111011101110111011101110111011101110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111010100100001000100010011011110000111011110000111011110000111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010000111011110001000100010000111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100010001000100010001000100010011001110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000010010001000010001000100010001001000100010001000100010001000100010000100010010001000100010000100100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101000011001100110011001100110011001100110011010001000011001101000101010101000100010000110011001101000011001100110011001100110010001101000100010001000100010001000100010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100001100110011001100110011001100110011001100110011001100110011001101000011010001000100010001000100001100110011001100110011001100110011001100110011001100110011010001000100010001000101010101010110011001100110011001100110011001100110011001100110011001010101011001100110011001010110011001010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101000100010101100101010101010100010001000101011001100110011001100110011101100111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101111000100001110111011101110111011110000111011101111000011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100001110111010100100001000100010010011110000111100010000111100010000111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010000111100010001000100001111000100010001000011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011001000010010000100010010010101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100100011001000110010000100010001000100010001000100010001001000010001000100010001000100010001000100010001000100010001001000010001001000010010001000100010001000100010001000010001000100010001000100010001001000100010001000100010001000100010000100010010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101010011001100100011001100110011001100110011001100110011010001000100010001000100001100110011010000110011001100110011001100110010001101000100010001000100010001000100001101000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100001100110011001100110011001100110011001100110011001100110011001101000100010001000100010101010110011001100110011001100110011001100110011001100110011001010101010101010110011001100101010101010101010101010101011001100110011001100110011001100110011001100110011001010110011101100110011001010101010101000100010101100110010101000100010001000101010101100110011101110110011001100111011101110111011101110111011101110111011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000100010001000011110001000100010001000100010001000100001111000100010001000100001111000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011000100001000100010010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001000010001000100010010010001110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000110010001000110011000100100010001000100001000100010001001000010001000100100001000100010001000100100001000100010010001000010001001000100010000100010001001000100001001000010001000100010001001000010001001000100010001000100010001000100001000100100010001000100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101000011001100100010001100110011001100110011001100110011010001000100010001000100001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010101010101010101100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101100110010101010101011001100110010101010101010101010110011001100110011001100101010101000100010101010101011001010100010001010101010001010110011001100110011001100111011101100110011101110111011101110111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101111000100001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011000100001000100010010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001000100001001000010001001101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010000100010010001000010010001000010010000100010001000100010010001000010001001000010001000100100010001000100010001000100010001000100010001000010001000100100010000100010010001000100010001000100010001000100010001000010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100010001100110011001100110011001100110011001100110100010001000100001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010101010101010001000101010101100110011001010110011001010101010101010101010101000101010101010101010101010101010101010101010101010110010101010101010101100110010101010101010101010110011001100110011001010101010101000101010101000101011001100101010101010100010001010110010101010101011001110111011001100110011001110111011101110111011101100110011001100110011001100111011101110111011101110110011101111000011101111000011001010101011001110111011101110111011101110111011110000111100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011000100001000100010010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000100001001000100001001001100111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100100010001000010001000100010001000100100010000100010010001000010010000100010010000100010010001000100010001000100010001000010001000100010010000100100001001000100010001000100010001000100001000100100010000100100010001000100010001000010001000100100010000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010101010101010001000100010101100110010101100101010101010101010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010110011001100110011001010101010101000101010101010101011001100110010101010100010101100101010101010110011001100110011001100110011001100110011101110111011101100110010101010101010101010110011101111000011101010101010101110111011101111000011001010101010101111000100010001000011101010101011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110001000100010001010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000100001001000010001001001010111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010001000100010001000100010010001000100010000100010010000100100010000100100010001000100010001000100001001000100001001000100010001000100010000100010010001000100010000100010001001000100010001000010010001000010001001000100010000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010101010100010001000100010101010101011001010101010101010100010001000100010001000100010101010101010101010101010101010101010101100101010101010101010101010110011001010101010101010101010101100110011001100110010101010101010101010110011001100110010101000100010101100101010101100110011001100110011001100111011001010110011001100110011101110110010101010101010101010110011101110111011001010100010101100111100010000111011001010101011110001000100010001000011001010101010101111000100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110001000100010001010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110110001000100001000100100001001001000111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100010010000100010001001000010010001000010010001000100010001000100001000100010001000100010010001000100010001000100010001000100010001000100010001000100001001000100010001000010010001000100010000100010010001000010010001000100010000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000011010001010100010001000100010001010100010001010101010101010100010001000100010001000100010001010101010101010101010101010101010101100110011001010101010101010110010101010101010101100101010101010110011001100110010101010101010101010110011001100110010101010100010101010101010101010101010101100110011001100110010101010101011001100101010101100110010101010101010101010111011101110110010101010101010101100110100010000111011101100110100010001000100010000111011001100101010101111000100001100101011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000001000100010001010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111001100100010001000100001001001000111011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010010000100100010001000100010000100010001001000010010001000100010000100100010001000100010001000100001000100100010001000100010001000100010001000100001000100010010001000100001001000100001000100010010001000010001001000100010000100010010001000100010000100010001001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100001100110100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110010101010100010101010101010101010101010101010110011001010101010101010101010101010101010101010101010101010110011001100110011001110110010101010101010101010101011001110110011001010110100010001000100010000111011101100101010101111000011101010101010101111000100010001000100001110111100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000001000100010001001110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111001100100010001000100010001000110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100100010001000010010000100010010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010000100010010001000100001000100100010000100100010001000100010001000010010001000100010001000010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010001010100010101010101010001000101010101010101010101010101010101010101010101010110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110010101010101010101010101011001110110010101010101011001111000100010000110011101100101010101010111011101100110010101101000100010001000100001010110011101010101100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010001000100010001001110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111011101110111011101110111010000100010000100100010001000100110011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100001000100010001000100010001001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010001000100100001001000010001000100100010000100100010000100100001000100100010001000100001000100010010001000100010000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010001010101010101010101010001000100010101010101010101010101010101010101010101010101010101010101010101010110011001100101010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011110000111011001010101010101100111011101110110011001101000100010001000011101100110010101000101011001010101010101010110011110001000100010000111011010001000011101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010000100010001001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001111000100001110111011101110111010100100010001000100010000100100101011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010010000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001001000100001001000100010000100100001001000100001001000100010001000100001000100100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100001101000100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010001010100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101010101010101010101010101010101011001110110010101010101010101100111011001100110010101110111100010001000100001100101010101010101010101010101010101010101011010000111011101110101010101100111011101100111011101110111011101111000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010000100100001001001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111010100100010001000010001001000100101011101110111011101110111011101110111011101110111011101110111,
	2400'b001000010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100100010001000100010001000100010000100010010001000100010001000100010001000100001001000010010000100100010001000100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011010001000100010001000100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010110010101100110011001100101011001110110011001100110011101110110010101010101010101010101010101010111011101100110011001100110011001100110011001100110011001100110011101100110011001100110011001100110011001100111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010000100010001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000011000100010001000010001000100100100011101110111011101110111011101110111011101110111011101110111,
	2400'b000100010001000100010001000100100001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100100010001000100010001000100010001000100010001000100010001000110011001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101010101010101010101010101010101010101010101010101100110010101010101011001010101010101100101010101010101011110000111011001010101011001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101111000100010001000011101111000100110001000100010001000100010001000100010001000100001110010000100010001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000010001001000100011011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010010001000100010001000100010001000100010001000100010001000100011001100100010001100110010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110100001100110011010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010000110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100101010101010101011001100101011001100101010101100110011101110110011001100110011101100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101111000100010001000100010001001100010001000100010001000100010001000100001110010000100100001000101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000010001000100010001000100010011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001100100010001100110010001000100010001000100010001000100010001000100010001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010000110100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001101000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101100101010101010101010101010101010101100101011001100110011001100110010101100101011001100110011101100110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101111000100010001000100010001000100010001001100010001000100110001000100101110010000100100001000101001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001000100010011010000111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110010001000100010001000100010001000100010001000110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010000110011010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001100110100010001000100010000110100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000101010001000100010001000100010001000100010001000100010001000101010101000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011110001000100010001000100010011001100110011000100110011001100101110010000100010001000100111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001000100010010110000111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001000110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000011001101000100010001000100010001000100010001000100010001000101010001000100010001000100010001000101010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101100111011101110111011101110111100001111000100010001000100110011001100110011001100101110010000100010010000100101000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100011001000100010001000100010010010000111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000110010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001100110011001100110100010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110100001101000011001100110011001100110011001100110011001100110100001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010001000100010001010110010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111100010011001100110011001100110000011000100010010000100101000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001000100010010001110111011110000111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100011001101000100010001000100010000110011001100110011001100110011001100110011001100110011001101000100010001000011001100100010001000110100010001000100010001000100010001000100010001000011001100110011001100100010001000100011001100110011001100110011001100110011001100110100001100110010001000110100010101000011001100110011001100110011001100110011010001000011010000110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010001010100010001010100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010000011000100010010000100100111100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100110011000100010011000100010001000100010001001100110001000100010001001100110011000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001000100010001101110111100010000111100001110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100011001100110011010001000100010000110011001100110011001100110011001100110011001100110011001101000110010000110011001100110010001000100011010001000100010001000100001100110011001100110011001100110011001000100010001000100010001100100010001100110011001100110011001100110011001100110010001000110100010001000011001100110100010001000011001100110100001101000011010000110011001100110011001100110011001101000100001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010100010001000100010001000100010101010110011101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010001000100100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000100010001001110111011110001000100010001000011110001000011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100010001001010101001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100011001100110011010001000100010000110011001100110011001100110011001100110011011001100010001001010110010000100010001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110010001101000100010001000100001100110011001100110010001101000011001100110011001100110100010101010100001100110011001100110011001100110011001100110100001100110011001100110011001100110011010001000100010001000101010101010101010101010100010001000100010001000100010101010101010101010101010101010101010001010101011001010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010010001000100101100010001000100010000111011110001000100001111000100010001000100010001000100001110111100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010000101001000100010001000100010001001101000100010001000100010001000100010001000100010001000,
	2400'b001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011010001000100001100110011001100110011001100110011001100110011011001100011001101000100010000110011001100110010001100100011001100110010001000110011001100110011010001000100010000110011001100110011010001000100010101010011001001000101010101010101010101010101011001010101010101100100001100110011001000100010001100110011010000110011001100110011001100100010001000110100001101000100010000110011001100110011010001010101010101100110011001100110011001100110011001010110011001100110011001100110011101110111011101110111010101111010101110100110011001100110011101110111011101100110011001100101010101010101010101010101010101010101011001100110011001110110011001010110010101100101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010011000100010000111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110011000100010010001000010101100010001000100010001000100010001000100010001000100010011001100110011000100110011001100110011000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000100010001000100010001001101001100110011001100110011001100110011001100110011001,
	2400'b010000110011001000010010001000100010000100100010001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100100011001100110011001100100010001100110011001100110100001100100011001100110010001000100011001100100010001000100011001100110100010001010101010101000100010001000100010101000100010001010100001100110100010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100001100110011010001000110011101110111011101110111011101110111011110000111011101100111011110001000100010001000100010001000100010001000010101101000100110011000100001110111100010000111100001110111011101110110011001100111011101110111011101110111011101110110011010001000011101101000100010001000100010001000100010001000100010001000100010001001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110001000100010001000100010001001101010011001100110011001100110011001100110011001100110011001100110001000100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010000100000100010010001000010100100010001000100010011001100110011001100110011001100110011001100110011010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110100111001000100010001000100010001001011010101010101001100110011001100110011001100110011001,
	2400'b010001000011001000010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100100010001100100010001000100010001000100011001100100010001000100010001000100010001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100001101000100001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001010111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001101000011110001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010000111011101111000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010111010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010011001100110011001100110001001100110010101000100010001000100010100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011000001000100010001000100010001001001001101010101010101010101010101010101001100110101010,
	2400'b001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010101010101010101100110011001100110011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010000111011110001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101110111010101010101001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010000111011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010000111011101111000100010001000100010011001100010001000100010001000100010011001100010011001101010101010101010101010101010101010101110110111000100010001001000010100101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100100010001000100010001000111001101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001000100010001000100011001100110011001100110011001101000011001101000011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110100010001000100010000110011001100110011001101000100010001000100010001000100010001000100010000110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101011001100110011001100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101101000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110101010100110011001101010101001100110011001100110011001100110011000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010011001100110011001100110011001100110011010101010011010101010101010101010101010101010101010101010101010101010111010100110101011101110111011101110111011101110111011101111001000001000010001001000010011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010000100010001000100010001000101000101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110100010000110011001100110011001100110011001100110010001100110011010001000100010001000011001100110011010000110100010100110010001000100011001100100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011010000110011001100110011001100110011001100110011001100110011010001000011001100110011001100110011010001000100010001000100010000110011001100110011001100110011001100110011010001000011010000110100001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001010100010001000100010001000100010001000101010101010110011001100110011001100111011101110111100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010011001100110011001100110011000100010001000100010001000100010001000100001110111011101110111011101111000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010111011101111001001001000010001001000010011101011001011101110111100101110111100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010100100010001000100010001000100110101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100100011001100100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000110010001000100011001100110011010001000100010000110011001100110011001100110010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110100001100110011001100110011001100110100001100110011010001000100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010001000100010101010100010101010101010101010101011001100110011001100111011101110111100010001000100010001000100010000111011101110111011101100110011001100110011001100110011001100110011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010000111011101111000100010001000100010001000100010001000100010001000100110011001101010101011110111011101110111001100101110111011101110111011101110111011101110111011101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100110011001011101111001100101110111011101110111011101110111011101111001010001000010001001000010010101011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000100010001000100010001000100101101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010101010101011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000100110011001100110001000100010001001100110011001100110011001100110011001100110011010101010101010101010101010101010101011101111001101111011111110111011011100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110111011101110111011110011001100110011001100110011001100101111001100101111001100110010111011101110111011101111001011001100010001001000010010100111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010011000100010001000100010001000100100101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000110011001100110011001100110010001000100010001000100010001000100010001100110011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001010101011001100110011001100111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101011101111001101111011111110111011101101110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100101110111011101111001100110011001100110010111100101111001011010000010001000100010010100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011100100010001000100010001000100011100010011001100110011001100110011010100110101010,
	2400'b001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101011001100110011001110110011001100110011001100101010101010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110101011101110111010101010101010101010111011101111001101111011111111111011101101110011001100101110111011101110111011110011001011101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001100101111001100110011001100101110111100110011001100101110111011110011001011101111001100110011001100110011001011010100010001000100010001011111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010100000100010001000100010001000100011100010011001100110011001100110101001100110011001,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000011001100110011001100110011001100110011010000110011010001000100010000110011001100110011001100110100010001000100010001010101010101010101010101010101010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001110111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001101010101011110011001011101010101010101010111011101111001101111011111111111011101101110011001100110011001011101110111011101110111010101111001100110011001100110010111011101110111011101110111011101110111011101110111010100110011010101110111011101110111011101110111011101110111011101110111100110011001100110011001100110010111011110011001100110011001100110011001011101111001100110011001100110011001100110011001100110011001100110011001100101110111100110010111011011000010001000100010001011011001100110011001100110011001100110011001100110011001011110010111011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001000010000100010010001000100010100010101010101010101010101010101010101010101010,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001000011001100110100001100110100010001000100010001000100010001000100001100110011001101000100010001000100010001010101010101010101010101010101010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101100110011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011110001000100001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101011101110111011101110101010101010111011101111001101111011111111111111101101110011001100110011001011101110111011101110111011101111001100110011001100110011001100110011001011101110111011101110111011101110111010101010101011101110111011101110111011101111001011101110111011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010111100110011001100110011001100110011001100110010111100011000010001000100010001010111001100110011001100110010111011110011001100110011001011110010111011101110111011101110111100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101001010010001000100010001000100010011110111011101110111011101110111011101110111011,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100001100110011001101000100010000110011010001000011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100101010101010101011001110111011110000111011110001000100010000111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001101010111011101010101010101010111011101110111011101110111010101010111011101111001101111011111111111111101101110011001100110011001100110011001011101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011110011001011101110111011101010101011101110111011101110111011101110111011101110111011100000010001000100010001010010111011101110111011101110011001101110111011101110111011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101001010010001000100010001000100010011010111011101110111011101110111011101110111011,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011001100110011001100110011001101000101010101000101010101000100010001010100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001110111011001100110011001100110011001110110011001100101011001111000100010001000100010001000100010001000100010001000100001110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011001100110001000100010011000100110011000100010001000100010001000100110101001100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011010101111001101101110101010101010111011101110111011101110111011101110111011110011001110111111111111111111101110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111010100110001010101110111011101010101001100110011001100110011001100110011001100110001001100110011001011100010001000100010001001110011010101010101001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101110101010101001100010000100100010001000100010010110111011101110111011101110111011101110111011,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100010001000011110001001101010101001100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001101010101010101010101010101010111011101110111011101110111011101110111011110011001110111111111111111111101110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101000011101111000100110101010101010101010101010101001100110011001100110011001100110011001100110011010100000100001000100010001001110101011101110111011101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110001000100110011001100110011001100110011001100110011001100110011001101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101010101010101010101010101001110010001000010010001000100010010110111011101110111011101110111011101110111011,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011001100110011010001000011001100110011001100110011001100110011001100110011001100110100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000011001101000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101000100010001010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110010101100110011101110111011101100111100010001000011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011010101010101010101010101010100110011000011110000111011101111000100110001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101010101010101010101010101110111011101110111011101110111011101111001110111011111111111111101110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100110011010101110111011101110111100110011001100101110111011101110111011101110111011101110111011101100110001000100010001001010011100110011001100110010111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011010101010101010100110001001100110101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111010101010101011101010101010101010000010001000100010001000100010010010101011101110111011101110111011101110111011,
	2400'b001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001101000011010000110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011101110111011101110111011101110111011101110111100010001000100010000111011101110111011101110111011101110111011110000111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110101010101010101010101010101010101010101011101110111010101010101000100010001000100010001000100010011001100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010111011101110111011101110111011101111001110111011111111111111111110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000001000100010001001010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001100110011001100110011001100110011001100110011001100110011010101010101001101010011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000011001000100010001000100010001110011011101110111011101110111011101110111011,
	2400'b001100110011001100110011001100110011001100110100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001110111011101110111011101110111011101111000100010000111011110001000100010000111011101110111011110001000011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000111100010001000100110101010101010011001100010001001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011110011011110111111111111111111111110110111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001010001000100010001001001111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101111001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101110111010101010011001100110011001100110011001100110011001101010011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110011001100110000100001000100001001000100010001110001010101010101010101010101010101010101010,
	2400'b010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010101010101010101010101010101000100010001000100010001000100010101010101010101010101010101100110011001100101010101010101010101100101010101010101010101010101010101010101010101100110011001100110011001100111011101110111011101110111011101110111011101111000011101110111100010001000100010001000100010001000011101110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101100110011101110111100010001001100110101010100110011000100010001000100010001001101010101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011110011011110111111111111111111111110110111001100101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001100001000100010001000101101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100101110111011101110111011101110111011101110111011101110111011101110111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100110011000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000100001001000100010001001111010101010101010101010101010101010101010,
	2400'b010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100101010101100101010101010101011001010101010101100101010101100101011001100110010101100110011001010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001011101010101010101010101011001100110011110001000100001110111011110001001100010101010101010111011101110111011101110111011101110111011101110111011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011011110111111111111111111111110110111001100110010111100101111001100110011001100110011001100110010111010100110011010101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001110001000100010001000101101100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010010111011110011010101010111011101110111011101110111011101110111011101110111011101010111010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100110000101001000100010001000010010001001101010100110011001100110011001100110011001,
	2400'b010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101100110011001100101011001100110010101010110010101010101010101100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010000111011101110111011001010101010101010101010101100101010101100110011001100110011101110111100010101011101110111011101110111010101010101010101110111010101010101011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101011101110111011101110111011101110111011110011001110111111111111111111101110110111001100101110111011110011001100110011001100110011001100101110010111011101111000011101111000100010001001100110011010100110001000101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010000001000100010001000101011011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100101110110011001100110100010101011101010101011101110101010101110101010101010011000100010011000011110001000100110101010101010101011101110111011101110111010101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101010101010101010101001100110011001100110011001100110011001100110011001100110011001100010000110001000010001001000100010001001011001100110011001100110011001100110011001,
	2400'b010101010101010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011001100110011001100110011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000011101110111011101110111011101110111011101110110011001100110010101100110011001111000100010001000100010001000100110011001100110101010101110111011101110111011101110111011101110111010101010101010101010101011101110101010101010101010101010101010101010101010101010101011101010111011101010111011101110111011101110111011101110111011101111001101111011111111111011101110110111001011101110111011101110111011101110111100110011001100101110000111011101111000100110011001100001110111011101110111100010001001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101111001011101111001011110010111100110011001100101111001100101111001100110011001100110011001100110011001100110011001100110011001100110011001100110010010010000100010001000101001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110101001011101100110011001100110011001111000100110011001100110001000100110011000100001110110011001100110011001100110011110001000100010011010100110011001100110000111011101110111011110011010101010101010101010101010101010101010101010101001100110011010101010011010101010101010101110111010101010101010101010101010101010101010101010101010101110101010101010111011101110111010101010111011101110101010101010101010100110011001100110011001100110011001100110010111001000100010001000010001001001011001100110011001100110011001100110011001,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110110011001100111011110001001100110011001100110011001100110011001100110011010101010101010101110111011101110111011101110111011101010101011101110111011101110101010101010101010101010101010101010101010101010101011101010101011101010111011101110111011101110111011101110111011101111001101111011101110110111011101110011001011101110111011101110111011101110111011101110111011101110010111011101110111100110011010100110001001100110011001101010111100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110011001100110011001100110011001100101111001011110010100010000100010001000100111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010010111011001100110011001100110011001100110011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100111011101100110011001100110011001100110011001111000100110101001100110001000100010001000100010001000100010001000100010001000100010011011110010111010101010101010101010101010101010101010101010101010101010101010101010101011101010001000100010011001101010111010101010101010101010101010101010101001101010011001100110010111001100100010001000100001001001001010101010101010101010101010101010101010,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111100010001000100010001000100010011000100010001000100110011001100110011001101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101011101010111011101110111011101110111011101111001100110111011101110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110011001100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110010100011000100010001000100111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010000111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001100110011001100110011001100110011001100110011001100110011001111001101010101010101010101010101010101010101010101001100110011001100010011000100010011000011101100111011101110111100010101011101010101010101010101010101010101001101010101001100110011000001100100001000100100010001000111001101010101010101010101010101010101010,
	2400'b010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100101011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001101010101010101010101010101010101010101010101001100110001000100001110111011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111100010011001100110101001100110011001100010001000100110011001100110011001100110101001100110011010101010101010101110111010101010111011101110111011110011001011101110101010101110111010101010101010101010101010101010101010101110111011101110111011101110111011101110111100110011001100110011001100110010111011101110111011101110111011101110111100110011001100110011001100110011001100110010111011101110111011101110111011101110111100110011001100110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110100000100010001000100101001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101001100110000111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101111000011101110111011101110111011101110111011101100110011101110110011001100110011001100110011101111000100010001000100010001000100110011001100110101001100110010111001100100001000100100010001000111000100110011001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110101010101010101010101010101001100110011000100010001000100010001000100001110111011101110111011101110111011101110111011101100110011001100110011001110111011101110111011101110111011101110111011110001000100010011001101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010111011101010101010101010101010101010101010101010101011101110111011101110111011101110111100110011001100110011001100110011001100110010111011101110111011110011001100110011001100110011001100110011001100110011001011101111001100110010111100110011001011110010111100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110100000100010001000100101001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010100110011001100010001000011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101100110011001010101011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111100010001000100010011000010000100001000100010001000100100111100110011001100110011001100110011001,
	2400'b011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001110111011101110111011101110111011101110111011101110111011110001000100110011001101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101110111011101110111011101110111011101110111011101110111100101110111011101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111100110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110101000100010001000100101000101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010011001100110011001100110001000011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011101110110010000100001000100010001000100100110100010001001100010001001100110011000,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011001110111011101110111011101110111011101110111011101110111011110001000100010001000100001110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101111000100010001000100010001000100010000111011110001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100110011001100110011010101010101010101010101010101010011001100110011001100110011000100010001001100110011001100110011001100110011001100110001001100110011001100110011001100110011001100110011011110011001100110010111010101010101011101110111011101110101010101010101010100110011001100110011001101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010100110000100010001000100010111101110111011101110111011101110111011101110111011101110101010101010101011101110111011101110111011101110111010101010101010101010101001100110011001100110001001100010011000100010000111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010110011001010101011001100110011001100110011001010101010101010101011001100101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100101011001100110010000100001000100010001000100100101011101110111011110001000100010001000,
	2400'b100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110101010101010101010101010101010101010101010101010101001100110011000100010001000100010001000100010001000100010001000100010001000100010011001100010001001100110011000100110011010101110111011101110101001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010011001100110011001100010001000100010000101000100010001000100010110101110101010101010101010101010011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110001000100010001000011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001000100010001000100100100011001100110011001100110011001100110,
	2400'b100010001000100010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110001000011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100110011010101010101010101010101010101010101010101010101010101010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011010101010011000100010001000100110011001100110011001100110011001100110011001100110001000100010001001100110011001100110011001100110011001101010101010101010101011101110101010101010101010101010101011101010101010101110111011101110111011101110111011101010111011101110101010101010101010101010101010101010101010101010101011101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010000110000100010001000100010101100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011001100110011001100110011000100010000111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001000100010001000100100100011001100110011001100110011001100110,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100010000111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001001100110011001100110011001101010101010101010101001100110011010100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100110011001100010001000100010001000100110011010101110101001100110011001100110011001100110011010101010011010101010011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101000001000010001000100010100100110011001100110011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010011001100110001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010000111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101100110010101010101010101100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000100001000100010001000100100011011001100110011001100110011001100110,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100001110111011101110111011101110111011001110110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100110011001101010101010101010101010100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001101010101000100010001000100010001000100010011000100010011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001000010001000100010011100110101010101010101010101010101010101010101010101010011001100110101010101010101010101010101010101010011001100110011001100010011001100110011010101010101010101010101010101010101001100110011001100110011001100110011001101010101001101010011001100010011001100110011001100110011001100110001000100010001000011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100001000100010001000100010011011001100110011001100110011001100110,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110000111100001110111011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100110011001101010101010101010101001100110011000100010001000100010011001100110001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101111000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100010001000100010011100110111010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010100110011001100110011001100110101010101010101010101010101010101010101001101010101010101010011001100110011001100110011000100010001000100010000111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110010101100110010101010110011001100101011001100110011001100110011001100111011101110110011101110111011001100110011001010101010101010101010101010101010101010101010101010101010101010101010100100001000100010001000100010011010101100110011001100110011001100110,
	2400'b011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010011001100110011000100010001000100010001000100010001000100010011001100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010001000100010001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010100110011001100110011001101010101010101010101010101010101010101010101010101010101001001100010001000100010010100010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001100110011001100110011001100010011000100110011001100110011001101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011101110111011101110111011001100110011001100101010100110001000100010001000100010010010101100110011001100110011001100110,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011110001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000100010011001100110011001100110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000100001111000100001110111011101111000100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011001010000010001000100010010011110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001100110011010101010011010101010011001100110011000100010001000100110011001100110011001100010001000100010001000100110011001100110011001100010001001100010011001100110101001100110011001100110011001100110011001100110011001100110011001100010000111011110001000100110011000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110001000011110001000011101110111011101110111011101110111011101111000011101111000100010001000100010001000100010001000100010001000100010001000011101110110011001100110011000110010000100010001000100010010011001100110011001100111011101110111,
	2400'b011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101111000100010001001100110101010101010101010100110001000100010001000100010001000100010001000100010001000100010001001101010101001100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001001100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001001100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000010000010001000100010001011010011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010011001100110011001100110011001100110011010101010101001100110001000011101110111011101110111011101110111011101110111011110001000100010001000100010011001100110011001100110011001100110011001100110101010100110011001100110011000100010001000100010001000100010001000100010001000100001111000101010101001100110001000100010000111100001110111011101110111011101110111011101000001000100010001000100010010011010001000100010001000100010001000,
	2400'b011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010000111100010001000100010001000011101110111011101110111011110000111011110001000100010001000100110101010101010111011101110111010100110011001100110011001100110011001100110011001100110011011110011011011101010011001100110011001100110011001100110011001100010001000100010000111011101110111011101110111011101111000100010011000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001001100110011001100110011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000010100010001000100010001010110011000100010001000100010000111011110001000100010000111100010001000011101111000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001001100110011001100110101010101010101001100110001000011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001001100110101001100110011001100110001000100010001000011101110111011101110111011101010010000100010001000100010001011010011000100010001000100010001000,
	2400'b011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011110001000100010001000100010001001100110011001100110011001100110011001100110001000100010000111011101110111011101100110011001100110011001100110011001100110011001100110011001100111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001110111011101110111011101110111100010000111100010001000100010001000100010001000100001110111011101110111011101110111100001111000100010001001100110101011101110111011101010101001100110011001100110011001100110011001100110011010101111001011101010101001100110011001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011001100010001000100010001000100010011001100010011000100010001001100110011001100110011001100110011001100110011001100110011000100010001000100010001000010100010001000100010001010010001000100010000111011110000111011101110111011101110111100010001000100001110111011101111000100001111000100010001000100010001000100010001000100010001000100010000111011110001000011101110111011101110111011110001000100010001000100010001000100001110111011101110111011101110111011101111000100010001000100010001000100010001000011101111000011101110111011101110111100001110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011010101010101001100110011001100110011000100010001000100010001000100010000111011101010010000100010001000100010001010110001000100010001000100010001000,
	2400'b011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100110001001100110011001100110011001100010001000100110001000100110011001100110011001100110011001100110001000100010001001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100001110111011101110110011001100110011001100110011001100110011101110111011110001001100110011001100110001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101111000100010001000100010001000100010000111011101110111011101110111011101110111011110000111011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011010110011011011101010011001100110011001100110011001100110011001100110011001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100010001000100010001000011000100001000100010001001101111000100001110111011101110111011101110111011101110111011101110111100010000111011101110111011101110111011110001000100010001000100010001000100010001000100010001000011110000111011101110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010001000100010000111100001100010000100010001000100010001010001110111011101110111011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011010101110111011101010011001100110011001100110011001100110011001100110011001100110001000100110001000100010001000011110001000011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100010011001100010001000100001111000011000100001000100010001001101111000100001110111011101110111011101110111011101110111011101110111100010000111011101110111011101110111011101110111011101110111011110001000100010001000100010001000011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101111000011110001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101100010000100010001000100010001001101110111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000111011101110111011110001000100010001000100001110111100001111000100010000111011101110111011101110111011101100110011001100101010101010101010101010110011001100110011101111001100110011001100110011001100110011001100110011001100110001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011001100110011000100010001000100010001000100110011001100110011001100110011001101110111010100110011001100110011000100010001000100010001000100010011001100110001000100010011001100110001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010001000100010001000100010001000100010001000011000100001000100010001001101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101100011000100010001000100010001001101100111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100110011001100110011001100110011001110110011001100110011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101011001111000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010001000011101110111011101100110011001100110011001100110011001110111011101110111011101110111011001110111011101110111011110000111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011010101111001011101010011001100110011001100110001000100010001000100010001000100110011001100110011001100110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011000100001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011000100010001000100010001001001100111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001010101011001100110011001100110011001100110011001110111011101110111011101110110011001100110011001010101010101010101010101010101010101010101010101100111100010001000100010001001100110011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110000111011001100110011001100110011001100110011001100110011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001001100110011001100010001000100010001000100010001000100010001000100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011110111011011101010101001100110011001100110011001100110011001100110001000100010011001100110011001100110011000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011110000111100001111000100010001000011101110111011101110111011110000111011110001000100010001000100010000111100001110111011101110111011000110001000100010001001001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011000100010001000100010001001001100111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101000100010101100110011001100110011001110111100010001000100010001000011101110111011101110111011001100110010101010101010101010101010101100110011110011001100110011001100110011001100110011001100110011001101010101010101010101010101010011001100110011001100110011000100010001000011101110110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001111000100010000111100001110111011101110111100010001000100001111000011101110111011101110110011001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101100111011101101110010111010101010101010100110011001100110011001100110011001100110011000100010011010101010101001100010001000100010001001100110011000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011100110001000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001100111011101110111011101100111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011000100010001000100010001001001010111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101000100010101100110011001100110011001100111011101110111011101110111011101110111011101110110011001100110010101010101010101010101010101010110011001111000100010011001101010101010101010011001100110011001100110011001100110011001101010101010101010011001100110000111011101110111011001100101010101010101010101100110011001100101011001100110011101100111011101110111011101110111011001111000100010001000100010001000100010001000100010001000011101110111011101110111011101110110011001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100010001000100010001000100110101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010111101111011101110110111001011101110111011101110111011101010101010101010101010101010101010100110011001100110101010100110011001100110011001100110011001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000001000100010001001001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110011001100110011001100110011001100111011101110111011001100111011001100110011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100000100010001000100010001001001010111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100110010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101000100010101100110011001100110011001100110011101110111011101110111011101100110011001100110011001100110011001100101010101010101010101100110011101111000100010001000100110011001101010101010101010101010100110011001100110011000100010011000100110011001100110011001100110011000100001110110011001010101011001100110011001100110011001100110011101110111011101110111011101110111011001101000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001110111011110001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011000100010011001100110011001101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101011101111001110111111111111111011011100101110111011101110111011101110111011110011001100110011001100101110111010101010011001100110011001100010011001100110011000100010011001100110001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101000001000100010001000101000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101110111011101100110011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001110110011001100111011001110111011001100110011001110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100000100010001000100010001000101010111011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010100010101100110011001100110011101110111011101110111011101110111011101110110011001100110011001100110011001100110010101010101010101100110011110001000100010001000100010011001100110011001100110101010100110011001100110011001100110011001100110011000100110011001100010001000100010000110011001010101010101100110011001100110011001100110011101110111011101110111011101110111011001111000100010001000100010001000100010001000100010001000100001110111011101110111011101110110011001110111100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010011001100110011001100110011001100110101010101010011001100110011001101010101010101010101010101010101010101010101001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010111101111011111111111011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011001100110011001100110011001100010011000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110110011101000001000100010001000101000111011101110111011101110111011101110111011101110111011101100110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100100000100010001000100010001000101000110011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101000100010101100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001110111100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001110111011110001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111101111111111111111011001011101110101010101010101010101010101010101010101010101010101001100110011010101010101010101010111011101110101010101010101010101010101010100110011001100110011001100110011001100110011001100110011000100010001000100010001000011101110111011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101100111011001100110011101110111011101110110011101010001000100010001000101000111011101110111011101110111011101110111011101110110011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011001100110011001100100001000010001000100010001000101000110011101110111011101110111,
	2400'b011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101000100010101100110011001100110011101110111011101111000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110011001100110011001100110011001100110011101110111011110001000100010000111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011101111000100010001000100010001000100010001001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101111001110111111111111111011011011101110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001001100110011001100110011001100110001000100010001000100110011001100110000111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100111011001100110011101110110011001100110011001100110011001100110011101010001000100010001000100110110011001110111011101110110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101100110011101110111011101100110011001100100000100010001000100010001000101000110011101110111011101110111,
	2400'b011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110010101010100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011001100110011000100010000111011101110111011101110111011101110111011101110111011101111000100010000111011101110111100010001000100001110111011001100110011001100110011001100110011001100110011110001000100010001000100010001000011110001001100110011001100110011001100110011001100110011001100110011001100110001000100001110110011110001000100010001000100010001000100010011001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101111001101111011111110111011001011101110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000100001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010001000100010001000100110110011101110110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011001100110011001100100001000010001001000100001000100110110011001110111011101110111,
	2400'b011101110111011101110111011110001000011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001110111010101010100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010110011101110110011001100110011001110111011101110111011101111000100010001000100010001000100010001000100010001000100110001001100110011001100110001000100001110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001110111011101100110011001100110011110001000100010001000100010001000011101111001100110011001100110011001100110011001100110011001100110011001100010001000100010000111011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101011101111001101111011111110111011011100101110111011101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011101110111011101110110011001100110011001100110011001100110011001100110011001010010000100010001000100110110011001100110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100100000100010001001000010001000100110110011001110111011001110111,
	2400'b011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101000100010101010110011001100110011001110111011110001000011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010000111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001110111011101100110011001110111100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101110111011101111001101111011111111111011011100101110111011101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001010010000100010001000100100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100110110011001110111011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001010101010101000101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001010100010101010101010101010101010101010101010101010101010101000100010101100110011001010110011001100110011101110111011110001000100001110111011101110111011101100110011001100111011001100110011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101111000100010001000100010001000100010001001100010001000100010000111011101110111011101110111011101110111011101110111100010011001101010101010101010101001100110011001100110011001100110011000100010001000100010001000100010011001100010001000100001110111011110001000100010001000100010001001100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101011101111001101111011111111111011011100101110111011101110101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010011001100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001010010000100010001000100100101011001100110011001100110011101100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100110110011001100111011101110111,
	2400'b011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101000101010101110111100010001000100010001000011101100110011001100110011001100110011001100111011101110111011101110111011101110111011101110110011001100110011001100110011001100111011101110111011101111000100010001000100010001000100010001000100110011001100110011001100110011010100110101010100110011001100110011001100110011000100010001001100110001000100110011001100110101010101010101011101110111010100110011001100110011001100110011001100110011001100110011000100010011000100010001000100010000111011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101111001101111011111111111011011100110010111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101010101010100110011000100010001000100010001000100010011001100010001000100010000111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010010000100010001000100100101011001100110011001100110011001100110011001010101010101010101010101100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100110110011001100110011101110111,
	2400'b011101110111011101110111011101110111011101110111011101110111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110011001010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010001000100010001111001100010011001100110011001100110011000100010001000011101110111011001100110011001100110011001100110011101110110011101100110011001100110011001100110011001100110011001100110011110001000100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010101010011001100110011001100110011001100110011001100110101011101110111010101010011001101010101001100110011001100110101001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111001101111011111111111011011100110010111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101110111010101010111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110001000100010000111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001010101011001010010000100010001000100010100010101010101010101010101010101100110010101010101010101010101010101010110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100110110011001100110011001110111,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110011001100101010101010101010101000100010001000100010001000100010001000100010001000100010101010101010101010100010001000101010101100110011001110111011110001000100010011001100110011001100110011000100010000111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111100010001000100010001001100110011001100110011001100110011001100110011001101010011010100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011010101010101010100110011001100110011001100110011001100110011001100110011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111010101010101010101111001101111011101110111011011100101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101010101010100110011001100110011001100110011001100110011001100110101001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100010000111100010000111011101110111011101110111011101110110011001100011000100010001000100010100011001100110011001100101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001010101010101010110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001010100010101010110011001100110010101100101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100100101011001100110011001100111,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000011101110111011101110111011001100110011001010101010101000100010001000100010001000100010101010101010101010101010101000101010101010101010101010101010101100110011001100111011101110111100010011001100110011001100110011000100010000111011101100110011001100101010101100110011001100110011001110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001001100110001001100010001000100010011000100110001000100010011001100110001001100110011001100110101001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101001100110011001100110011001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101011101110111011101010101010101111001101111011101110110111001011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101010101110101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000100010100100001110111011101110111011101100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000101010101000101011001010101010101010101010101010110010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100100101011001100110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001111000100010001000100010000111100010001000011101111000011101110111011101110111011101110111011101100110011001100110010101010101010101010101010101010100010101000100010101010101010101010110011001010101010101010101010101100110011001100110011001110111100010001001100110011001100010001000011101110110011001100110011001100110011001110111100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100010001000100110011001100110011001100110011001101010101010101010101010101010011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101111001101111011101110111011001100101110111011101110101011101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110001000100010001000100010001000100010001000100010001000100010001001100110011000100001110111011101110111011101110111011101110111011101110111011101110100000100010001000100010100100010001000100010001000100001110111011101110111011101100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101000101010101010101010001000100010101010101010101010101010101010101010101010100010101010101010101010101010101010101010101010101010101010101010101010100010001010100010001010101010101010110010101010101010101010101010101010110010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100000100010001000100010001000100100101011001100110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000011101111000100001111000011101110111011101110111011101110111011101110111011101110110011001100110010101010101010101100101010101010101010101010101011001100110011001100110011001010101010101010101010101010101010101100110011001110111011101110111011101110111011001110111011101110111011101110111011101111000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001001100110001000100010001000100010001000100110001000100010001001100110011001100110101010101010101010101010011001100110011001100110011001100110011010101010101010101010111011101110111010101010101010101010101001101010011001100110011001100110011001100110101001100110101010101010011001100110011001100110011001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111001110111011111111111011011100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010100110011010100110011001100110011001100110011001101010101010101010111011101110111011101110101010101010011001100110011001100010001000100010001000100110001001100110011001101010011001100110011001100010001000100001110111011101110111011101110111011110000101000100010001000100010100011110001000100010000111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101000100010101010100010101010101010001010101010101010101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010001010101010101010101010101010101010101010100010001000100010001000101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010100001000010001000100010001000100100101011001100110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011101111000100001110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101010101010100010001010101010101010101010101100110010101010101010101010101010101010101010101010101010101010110010101100110011001110111011101110111100010001000011101110111011101110111011101111000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010111011101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010101001101010011001100110011001100110011010100110101010101010101010101010101010101010011001100110101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111100110011001101111011111111111011011100110011001011101110111011101110111011101110111010101110111011101110111011101010111011101010101011101010101010101010101010101010101010101010101010100110101010101010101001101010101010101010101010101010101010101010101011101110111011101110111011101110101010100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010011001100110011001100010001000100010001000100010000110001000010001000100010011011101110111011001100110011001100110011001100110011001100110011001100110011001100101010101010101011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001010101010101010101010101010101010101010101010101010100010001000101010001000101010101000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100101010101010101010101010100001000010001000100010001000100100101011001100110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110110011001100101010001000100010001010100010101010101010101010101010101010110010101010101010101010101010101010100010001010101010101010101011001110111011101110111100010001000100001110111011101110111011101110111011110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101110101011101110011001100110011001100110011001100110001000100010001000100010011010100110011001100110011001100110011001100110011001101010011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010111011101110111011101110111011110011001101111011111111111011011100110010111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101010101010101010101010101010101011101110111011101110101010101010101010101010101010101010101010101010011001100110011001100110011000100010010111001000010001000100010010011110000111011101110111011101100111011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000101010101000100010001000100010001000100010001000100010001000100010001000101010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001010101010101010101010101010100001000010001000100010001000100100101011001100110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111010101010101010101010101010101010101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011101110111011101111000100010001000100010001000011101110111011101110111100010001000100010001000100010011000100010001000100010001000011101110111011101110111011101110111011110000111011101111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001001100110001000100010001000100010011001100110001000100010001000100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101110111011101110111011101111001110111111111111111011011100110010111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110011001100110011001100110011001100110011001100010001000100010001000100010000111001000010001000100010010011001110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100001000010001000100010001000100100101011001010110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001100110011001010101010101000100010101010101010101000101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100111011101110111100010001000100010001000100010001000100010000111011110001000100010001000100010011001100110011001100110011000100010001000011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001101010011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101001100110011001100110011001100110011001100110011001101010101010101010101001100110011010101010011001100110011001101010101011101110111011101110111011101111001101111111111111111011011100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101010101010101010011001100110101010101010101010100110011001100110011001100110001000100110011001100110011001100010001000100010000111001000010001000100010010011010001000100010000111011110001000100010001000100010011001100110011001100010001000100001110111011101110111011101100110011001100110011001010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101011001100101010101010101010001000100010001000100010001000100010101010101010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000100010001000100010001000100100100010101010101011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110011001100101010101010101010101010101010101010101010101010100010001000101010101010101010101010101010101010110011001100110011001100110011001100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011000100010000111011101110111011101111000100010001000100010001000100010001000100010001000100001110111100001111000100010001000100001110111011101110111011110001000100010000111011110001000100010001000100010001000100010001001100110011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101111001101111011111111111011101100110010111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010101010101010101010101010101010100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100010001000100010001011010011001100110011001100110011010101010101010101010101010101010101010101010101001100110011001100110001000100010001000100010000111011101110111011101100110011001100110011001100110010101010101011001010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100101011001010101011001100110010101010101010101010100010001000100010001000100010001000100010001010100010101010100010101010101010101010101010101010101010101010101010001000101010101010100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000100010001000100010001000100100100010101010101010101100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111100010001000100010001000100010001000100010001000100010001000100010000111011101110111011001100101011001010101010101010101010101000101010001000100010001000100010001010101010101010110011001100110011001100110011001100111011101100111011101110111011101110111011101111000100010001000100010001000100010000111011101110111011110001000100010011001101010101001100110011000100010001000011101110111100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010011010100110001000100010011001100010001000100010001000100110011000100110011001100110011001100110011010101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011110011001100110011001100110011011110111011111110111011011100101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010000010001000100010001011010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110001000100010001000100010000111011101110111011101100110011101100110011001100110011101110111011001110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000100010001000100010001000100100100010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110011001010101010101000101010001000100010001000100010001000101010101010101010101010101010101010110011001100110011001110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000011110001000100010001001100110101010101010101010101010011001100010001000100010001000100001110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010011010100110001000100010001000100010001000100010001000100010001001100110001000100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101111001100110011001100110011011110111111111111111011011100101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110001000100010001000100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101001100110101010010000010001000100010001010110011001101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011000011101110111011101110111011101110111011101100111011101110111011101110111011101111000100010001000100010000111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010011000100010001000100010001000100010100010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011001100101010101010101010101000100010101000100010001000101010101010101010101010101010101100110011001110110011001110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100110101010101110111011101110111011101110101010101010011001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001001100110000111100010001000100010001000011110001000100010001000100110001000100010001001100110011001100110011001100110011010101010101010101010101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011110011001101111011111111111111011100101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001010100010001000100010001010110101010101010101010101010101010100110011001100110011001100110011001100010001000100010001000100010011001100110011001101010101010101010101001100110011000100010001000100010000111011101110111011101100110011101110111011101110111011101111000011101110111011101110111011001100110011101100111011101110111011101110111011101100110011001100111011101110111011101110110011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010011000100010001000100010001000100010100010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010000111100010001000011110001000011101110111011101110111011101110111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100101010101010101010101010100010001000100010001000100010101010101010101010110011001100110011001100110011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100110101011101110111011101110111100110010111100101110101010101010101001100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100001110111011101111000100010001000100010001000100010001000100110011000100010001000100010001001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101011101110111011101110111011101110111011101111001101111011111111111111101100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000010001000100010001010110101010101010101010101010011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101100101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010001000100010101010011000100010001000100010001000100010011010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011110001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000011101111000100010001000011110001000100010000111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001010101010001000101010001000100010001000101010101000101010101010101011001100110011001100111011001110111011101110111011101110111011101110111100010001000100010001000100010001001100110101001100110101010101010111011101111001100110011001100110011001100110010111011101110111010100110011000011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101011101110111011101110111011101110111011110011001110111011101110111011011100110011001011101110111011101110111100110011001100101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010011100100001000100010001010010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100110011001100110101010101010101010101010101001100110001000011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100101010101010101010101010101010101100101010001000101010101010011000100010001000100010001000100010011010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110000111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110010101010101010001000100010001010101010101000101011101100101011001010101010101100110011001100110011101110111011101110111011101110111011101111000100010001000100010001001101010101010100110101001100110101010101010101010101110111011101111001011110011001100110011001100110011001011101010101001100110001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011110001000100001111000100010001000100010001000100010001000100010001000100110011000100010001000100010011001100110011001100110101010101010101010101010101001100110011001100110011010101010101010101010101010101010101011101110111011101110111011110011011110111111111110111011011100110011001011110010111011101110111011110011001100110011001011101110111011101110111011101110101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000100001000100010001010010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010011001100110011010101010101010101010101010101010011000011110000111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010110011001100110011001100110011110000111100010000111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010101000101010101010011000100010001000100010001000100010011010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111100001110111011101111000100010000111011101110111100010001000100010001000100001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110010101010101010101010101010101010101011110000110010101100110011001100110011001100110011001100110011101110111011101110111011101111000100001111000100010001000100110011001101010101010101010101010101010011001100110101001101010101010101010101011101110111011110011001100110011001100110011001011101110111011101110111011101110111011110011001100110010111011101010011000011101110111011101110111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000100110011001100110011010100110001001100110011001100110011001100110101010101010101010101010101010101110111011101110111011110011001110111011101101110111001011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000100001000100010001001110011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011000100010001000100010001000100010001000100110011001100110011001100110011000100010001000100010000111011101110111011110001000100010001000100010001000100010001000100001110111011101110111011001100110011001100110011001100110011001100110011001110111011101110111011101110110011101110111011101110111011101100110011001010101010101010101010101000100010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010001000100010011010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011110001000100010001000100001110111011101110111011110001000011110000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100101010101010101010101010101010001010101010101100110011001110111011001100110011001100110011001110111011101110111011101110111011101110111100010001001100110011001100110101010101010101010101010101010100110011001100110011001100110011001100110011010101010101010101110111011101110101010100110011001100110101010101010101011101111001100110011001011100110001000011101110111011101110111011110001000011110001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100010001000100010001000100110011001100110011010101010101001100110011001101010101010101010111011101111001101110111011100110010111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101001100110101010100100110001000100010001001010001010100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110101010101010111011101010101010101010011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010011001100110001000100110011001100110011001100110011001100110011001100110011001100110011000100001110111011101100110011001110111011110001000100010001000100010001000100001110111011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010001000100010011010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110011001100110010101010101010101010101010101100110011001100110011001100101010101100110011001100110011001100110011101110111011101111000100010001000100010001001100110011010101010101010101010101010101010101010100110011001100110001001100110011000100110001001100110011001100110011001100110011001100110011001100110011001101010101010101010101001100010001000011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010001000100010001000100010011001100110011010101010011001100110011001100110011001100110101010101010111100110111011101110011001011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100100110001000100010001001010001010101010101010101010101010101010101010101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010011001100110011001101010011001100110011001100110011001100110011001100110011000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110001000011101110111011001100101010101010101010101010101010101100110011001110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001100110011001100101010101010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010001000100100011010101010101010101010101,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110010101010101010101010101011001100110011001010101010101100110011001100110011001100110011001100110011001100111011101110111011101111000100010001001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010011001100110001000100010000111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001101010101011110011011101110011001100101110111011101110111010101010101010101010111011101010101010101010101010101010101010101010101010101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010100110011001100110011001100110011001100110101010100101000001000100010001001010001011101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100001110111011101110111011101110111011101110111011101110110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000101010001010011000100010001000100100001000100100011010001010101010101010100,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011001100110011001100101010101010101010101010110011001100110011001100110011101110111011001100111011001100110011101110111011101110111100010001000100010011001100110011010101010101010101110111011101110111011101110111011101110111010101010101001100110011001100110011001100110011001100110011001101010101010101010101011101110111100101110111011101010101001100110001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011010101010101010101110111011101110111011101110111011101010101011101110111010101010101010101010101011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101011101010101011101110101010101010101010101010101010101010101010101001000001000100010001001010001011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011110001000011101110111011101111000100001110111011101110111011101110111100010001000100010001000100010001000011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010001000100010001000100010001000100010001010101010101010011000100010001000100100010000100010011010001010101010101010100,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101111000100010000111011110001000100010001000100110011001100110101010101010111011101110111011101110101010101010101010101010101010101010101010100110011001100110011001100110001000100010001000100110011010101110111011101110111011101110111011101010101001100110001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110101010101010101010101110101010101010101010101010101010101110111011101110111010101010101010101110111011101110111011101110111010101010101010101010011001100110101010101010101010101010101010101010101010101110101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101101010001000100010001000101111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010011000100010001000100010001000100100010010101100110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011110001000100010001001100110011001100110011010101010101010101010101010101010101001100110011010101010101010101010101010101010011001100110011000100010001000100001111000100010001000100110101010101010101011101110111011101110111010101010011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101010101010101010101011101110111011101110111011101110111011101110111011101110111011101101100001000100010001000101101011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100010001000100010001001000010010011001110110011001100110,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001110111011101110111011110001000100010011001100110011010101010101010101010101001101010101001100110011010101010101010101010101010101010101010101010101010100110011001100110011000100010001000100010000111011110001000100010001001100110011001100110101010101010101001100110011001100110001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001101010011010101010101010100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101101100001000100010001000101011011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011101110111011101110111011101110111011101110100000100010001000100010001000100010010011001110111011001100110,
	2400'b011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011101111000011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011001100110011001100111011101110111011101110111011101110111011110001000100010011001100110101011101110111010101010101010101010101010101010101011101110111010101010101010101010101010100110011001100110011001100110011001100110001000100010001000100001110111011101110111011101110111100010001000100010001000100010001001100010001000011110001000011101110111100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001101010101010100110011010100110011001100110011001100110011001100110011010101010101010101010101010101010111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010101011101110111010101101100001000100010001000101001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010000111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110100000100010001000100010001000100010010011001110111011101110111,
	2400'b011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010011011101110111011101110111011101010101010101010111011101110111011101110111011101110111010101010101010101010101010101010101010101010101001100110011001100110011001100110011000100010001000100010001000100010001000100010011000100010000111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101110111011101110111010101101110001000100010001000100111001101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101001100110011001100110011001100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010000111011101110111011101110111011101100111011101100110011001100110011001100111011101110111011101110111100010001000100001110111011101110111011101110111011110001000100010001000100010001000100010000111011101110111011101110111011101110100000100010001000100010001000100010010011001110111011101110110,
	2400'b011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010011011101110111011101110101010100110011001101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110001000011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101110111010101110111011101110111011101110101001100110011001100110011001101010101010101110111010101101110010000100010001000100111001101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110100000100010001000100010001000100100010011001110111011101110111,
	2400'b010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010101110111011101110111010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110001000100010001000100010001000100010001000100010001000100110011001100110011010101010101010101010101010100110011001100110011001100110011001100110011010101010101010101010101010101010101001100110011001100110011001100110011001100110011010101010101011101110111011101110111011101110111010101010011001100110011001100110011001100110011001100110101010101110000001000100010001000100101001101010101010101010101010101010101010101010101001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100110011001100110011001100110001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100100001000100100010001000100010011001110111011101110110,
	2400'b011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100110011011101110111011101110111010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010100110011000100010001000100001110111100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100110011010101110111010101010101001100110011001100010001000100010001000100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101110111011101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110000010000100010001000100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000011101110111100010000111011101111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100000100100001000100100010001000100010011001110111011101110110,
	2400'b011001100110011001100110011001100111011101110111011101100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010011001100110101011101110111011101110111011101110111011101110111011101110111011101110111100110011001011110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101001100110001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001101010101001100110011001100010001001100010001000100010001000100010011001100110011001100010001000100010001000100010001000100010001000100010011001100110011001100110011010101110111010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100101110010000100010001000100010111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101001100110011010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100110011010101010101010100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010001000100010001000100010001000100010000100001000100001000100100010001000100010011001110111011101110111,
	2400'b011001100110011001100110011001100110011101110111011101100110011001100100010000110011010001010101010101010101010101010101010101010101010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110101010101110111011101110111011101110111011101110111011101110111011101111001100101110111011110011001100110011001100110011001011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010100110011001100110011000100110011010100110011000100010001000100001110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011000100010011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001101010101001100110101010101010101010101010101001100110011001100110011001100110011001100110011001100110000010000100010001000100010111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110101010101010011010101010101010101010101010101010101010101110111011101110111011101110111010101010101010101010101010101010101001100110011001100110011000100010011001100010011001100110001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010000100001000100001000100010001001000100010011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100101010101000100001100110100010101100110010101100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011000100010011001101010101010101010101010101010101001100110011001100110011001100110011001100110010011000100010001000100010110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010111011101110111011101110111011101110111011101010101010101010101010101010101001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100001000100010010001000100011011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110010101010101010101000100010001010101010101010101011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101010111011101110111011101110111011101111001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110001000100010001000100010000111011110001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110101010101010101010101010011001100010011001100110011001100110011001100110010011000100010001000100010101101010101001101010101010101010101001100110011001100110011001100110011001101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001110111011110001000100010000100001000010001000100010010001000100011011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110010101010110010101010110010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100010000111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110001000100010001000100010001000100110011001100110010011000100010001000100010100100110011001100110011001100110011001100110001000100010001000100010001001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111010101010101010101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010000100001000100001000100010010001000100011011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100001110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000011000100010010001000010100100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010011001100110011010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010111011101010101010100110011001100110011001100010001001100110001000100010001000100010000111011101110111011101110111011101110111011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010000100001000100001000100010010000100100011011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011101110110011001110111011001100110011101100110011001100110011001100110011001100110011001100110011001110110011001100111011101100110011001100110011001100110011001100110010101010101011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010011000011101110111011101110111100010001000011101110111011101110111011101110111011101110111100010001000011110000111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100110011010101010101010101010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100000100010001000100010011100010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100110011001100110101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100010001000100010001000100001110111011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010000100001000100001000100100010001000100011011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001110111011001110111011101100110011001100110011001100110011001100110011001100110011001110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010011001100110001000011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001001101010011001100110101010101010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101000100010001000100010011100010001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110000100001000010001000100100010001000100011011001110111011101110111,
	2400'b011101110111011101110111011001100110011001100110011001100110011001110111011001110110011101100111011101110111011001110111011001100110010101010101011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101001100110011001100110011001100110011001100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111100010011001100001110111100010011010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110000100010001000100010010011110001000100010011001100110001000100010001000100010001000100001110111011101111000100010001000100010001000100010011001100110101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001001100110011001100110011001100110011001101010011001100110011001100110011010101010011001101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100100010001000100011011110001000011101110111,
	2400'b011001110111011101110111011101110110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001110111011101110111011101110111011101110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011101010101010101010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010011001100110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101110111011110001001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101000100010001000100010010011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010011001100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100100010001000100011011110001000011101110111,
	2400'b011101110111011101110111011101110110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110110011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010111011101110111011101110111011101110111011101110111011101110101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110000100010001000100010010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001001100110001000100010011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100100010001000100011011110001000011101110111,
	2400'b011101100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011110001000011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010000110000100010001000100010001011010000111100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100010010001000100011011110001000100010001000,
	2400'b011001100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011000100010001000100010001000100010001000011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011110000111011101110111011110000101000100010001000100010001010101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100010001000100100011011110001000100010001000,
	2400'b011001100110011001100110011001100101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011000100010000111100010001000100010001001100110001000011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010000110000100010001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110101001100110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010000011000100010001000100010001000100100011011110001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101110111011101110101011101110101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001000100010011001100110001000011110001000100001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101000100010001000100010001010001110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010011000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010000011000100010001000100010001000100100011100010001000100010001000,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101000100010001000101010101000011010001000100010001000100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001110111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100110001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000011101111000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001000100010001010100010001010100010001000100010001000100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100001110111011101111000100010001000011101110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111100010001000011101111000100010001000100001110111011101110111011101110111100001110111011110001000100010001000100010011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100101010101010101010001000100010000110011010001000100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100001111000100001110111100010001000100001111000100010000111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011101111000011101111000011101110111011101110111100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010000111011101111000100010001000100010000111011110001000100010001000100010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101010101010101010001000100010000110011010001000100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011101110111011101111000100010000111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101111000100010000111100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101010101010101010101010101000100010001000011001101000100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110100010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110010101010100010001010101010001000100010001000100001101000100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010011001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100101010001000100010001000100010001000100001100110100010001010110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001101010111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010100010001000100010001000100010000110100010001010110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001100110100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001010101011001100101010001000100010001000100010000110011010001010111011001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001100110011001100110011001100110011001101100111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101010101000100010000110011010000110011010001010110010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010000110011001100110011001100110011001100110101011101110111011101100110011001110111011101110111011101110111011101110111011101110111011001010101010101010101010101010101010000110011001101000011001101000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100010001001100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010001000100001100110011001100110011001100110011010001110111011101100110011001110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101010000110011001100110011001101000100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011110001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010001000100010001000011001100110011001100110011001101000110011101100101010101100111011101110111011101110111011101110111011101110111011001100101010101010100010001010100010001000011001100110011001101000100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101000100010001000100001100110011001100110011001100110011010101100100010101010110011101110111011101110111011101110110011101100110011001100110011001010101010001000100010001000100001100110011001101000100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001010101010101000100010001000011001100110011001100110011001101000100010001010101011001100111011101110111011101110110011001100110011001100110011001010101010001000100010000110100010000110011001101000100010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101010101000100010001000100001100110011001100110011001100110100010001000100010101010110011101110110011101100110011001100110011001010101010101100101010101000100010000110011010000110011001100110100010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101111000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100101010101010101010001000100010000110011001100110011001100110011001101000100010001010110011101110110011101110110011001100101010101010101010101010101010101000100010000110011001100110011001100110100010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101010001010100010101010101010001000011001100110011001100110011001100110100010001010100011001100111011101110110011001100101010101010100010101010101010101010100010000110011001100110011001100110100010001010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101000101010001000101011001100110010101010101010001000011001100110011001100110011010001010100010101010110011001100110011001100101010101010101010001000100010001010101010000110011001100110011001100110011010001010101011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010000111011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010101010101010101010101010100010001000100010001000011001100110011001100110011001101000100010001000101011001100110011001100110010101000100010001000100010001000100010101000011001100110011010000110011010001000101011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101110111011101111000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101000100010001010100001100110011001100110011001100110011001100110011001100110011001100110100001101000101010101100110011001100110011001010101010001000100010001000100010001010011001100110011001100110011001101000101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010001000100010001000100010001000100010001000011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b010101010110011001100101010001000011001100110011001100110011001100110011001100110011001100110011010001000100010101010110011001100110011001010101010101000011001100110011010001000100001100110011001100110011001101000101010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101111000100001110111011101110111011110001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101100101010101010101010000110011001100100010001100110011001100110011001100110011001100110100010001000101010101100101011001100101010101010101010000110011001100110011010000110011001100110011001001000100010101010110010101100111011101100111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010000111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110011001010100010001000101010101010100001100100010001000100010001100110011001100110011001100110011010001000100010101010101010101010110010101000100010000110011001100110011001101000100001100110011001000110100010001010101011001100111011101110111011101110111011101110111011101110111011101100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010000111100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001010101010101010101010001000101010101010100010000110010001000100010001100110011001100110011001100110011001101000100010001000100010101010101010101010100010001000100001100100011001100110100001100110011001000110100010101010101011001100110011101110111011101110111011101110111011101110111011001010101010101010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110010101010101010001000100010001000101010001000011001100100010001000110011001100110011001000110011001100110011010000110100010001000100010001000100010000110100010000100010001100110011001100110011001000110100010101010101010101100110011101110111011101110111011101110111011101110110010101000100010001000100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110010101010110010101010101010101000100010001000011001100110010001000100011001100110011001100110011001100110011001100110011001101000100010001000100010000110011001100110010001000110011001100110010001000110100010101010101010101010110011101110111011101110111011101110111011001100101001100110011001101000110011001100110011101110111011101110111011101110111011101110111011101110111011001100110011001110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110010101010101010101010101010101010101010101010100001100110011001000100010001100110011001100110011001100110011001100110011001101000100010001000100001100110011001100110100001000100011001100100010001000110100010101000101010101010110011001110111011101110111011101110110011001010100001100110011010001000100010001000101010101100110011001110111011101110111011101110111011101110101010101100111011101100101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100110010101010100010001000101010001000011001100110011001000100010001000110011001100110010001100110011001100110011001100110100010001000011010000110011001100110011001100100010001100100010001000110100010101000100010001100110011101110111011101100111011001100101010001000011001100110011010001000100010001000101010101010101010101100110011101110111011101110111011001010101011001110110010101010110011001110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001101010111011101110111011101110101010100110011001100110011001100110011001100110011000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110010101010110011001100110010101000011001100110011001100110010001000100010001000100011001100110010001000110011010000110011001100110011010001000100001100110011001100110011001100110011001100100010001000110100010001000100010101010101011001110111011001100110010101000100010000110011001101000100010001000100010001000101010001010101010101010101011001100110011001110101010001010111011001010101011001100110010101010101010001000100010001000101010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011000100010011001101010111100110111011101110111011101110111011100101110101001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011001100110011001100101010101010101010001000011001100110011001100110011001000100010000100100011001100110011001000100011001100110011001100110011001101000100001100110011001100100010001100110011001000100010001000110100010001000100010101000101010101100110010101100100010000110011001100110011010001000100010001000100010001000100010001010101010101010101010101010101010101000011010101100100010000110100010001000100001101000100010001000100010001000100010001000100010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011011110011011101110111011101110111011101110111011101110111001011100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101100110011001100110010101100101010101000100001100110010001000100011001100100010001000100010001100110011001100100011001100110011001100110011001100110100010000110011001100100010001100110011001100100010001000110011010000110100001100110101010101100101010101000011001100110011001100110100010001000100010001000100010001000100010101010101010101010101010101010100001100110011010000110011001100110011001101000100010001000100010001000100010001000100010001000100010101010101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001101011001101110111011101110111011101110111011101110111011101110111011101101110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101100110011001100110010101010101010000110011001000100010001000100010001000100010001100110011001100110010001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000110011010001000100001100110100010101010100010000110011001100110011010001000100010001000100010101010101010101010101010101010101010101010101010000110010001100110011001100110011001101000100010000110100010001010101010001010101010001010100010001000100010001000101010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011010110011011101110111011101110111011101110111011101110111011101110111011101110110111001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b011101110111011101100110011001100101010101010100010001000100001100110010001000100010001000100010001100110011001100110011001000110011001100110011001100110011001100110011001100100010001000100011001100110010001000110011010000110011001100110011010001000100001100110011001100110100001100110011010001000100010001010101010101010101010101010101010101000011001000100010001000110011001100110100010001000101010101010100001101000101010101010100010101100110011001010100010001000100010001010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110101100110111011101110111011101110111011101110111011101110111011101110111011101110111011011100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111,
	2400'b010101110110011001100110011001100101010101010101010001000100010000110011001000100010000100100010001000110011001100110011001100110010001000110011001100110011001100110010001100100010001000100010001000110010001000110011001100110011001100110011001101000011001100110011001100110011001101000100010001000100010001010100010001000101010101010100001100100010001000100010001000100011001100110100010001000100010001000101010001000100010101010100010001100110011101110110010101010100010001000100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100111001101111011011101110111011101110111011101110111011101110111011101110111011101110111011100101010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001001000110011001100110011001010101010101010101010101000100010001000011001000100010001000100001000100100010001100110011001100110011001000100010001100100011001100100010001000100010001000100010001000100010001000100011001100100010001100110011001100110011001100110011001100110011010001000100010001000100010001010101010001010100010000110010001000100010001000100010001000110011001100110011010001000100010101000100010101000100010001010101010001010110011101110111011101100101010101000100010001000100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001101111011110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100011010101100110011001100101010101010101010101010100010001000100001100110010001000100001000100010010001100110011001100110011001100100010001000110011001000100010001000100010001000100010001000100010001000100011001100100010001100110011001100110011001100110011001100110011010001000100010001000100010001010101010101000011001000100010001000100010001000100011001100110011001100110011001101000100010101010101010101010100010001000101010101010101011001110111011101110110010101010101010001000100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010110111101101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110110,
	2400'b001000100010001001000101011001010101010101010101010101010101010001000100001100110011001000100001001000010001001000100011001100110011001100110011001000100011001100100010001000100010001000100010001000100010001000100011001000100010001000100011001100110011001100110011001100110011010001000100010001000101010101010101010000110010001000100010001000100011001100110011001101000100001100110011001100110100010001000101010101010101010001000100010101010101010101100111011101110111011101100101010101000100010001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011011111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110111001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110,
	2400'b001000100010001000100011010001010110011001010101010101010100010001000100010000110011001000100010000100010001000100100010001000100011001100110011001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100011001100110010001100110011001100110011010001000100010001000100010001000100001100100010001000100010001000110011001100110011001100110100010001000100001100110100010001000101010101100101010101000100010101100101010001010111011101110111011101110101010101000100010001000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110101101111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011101110111001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111,
	2400'b001000100010001000100010001000110100010101010101010101000100010001000100010000110011001000100010000100010001000100100010001000100010001100110011001000100010001000100010001000100010001000100010001000010010001000100010001000110011001000100010001100110010001000110011001100110011001101000100010001000100010001000011001000100010001000110011001100110011001100110011001100110011010001000100010001000100010001000100010101100110010101010100010101100110010101010110011101110111011101110111011001000100010001000100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110101101111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011101110111011010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111,
	2400'b001100100010001000100010001000100010001101000101010101000100010001000100001100110011001000100010001000010001001000010010001000100011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001100110011001100110011001100110100010001000100010000110010001000100011001100110011001100110011001100110011001100110011001101000101010101000100010001000100010101010110010101010100010001010110011001010101011001110111011101110111011101100100010101000100010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100110111110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011101110111011010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110,
	2400'b001100110010001000100010001000100010001000110011001101000100010001000100010001000100001100100010001000010001000100010001001000100010001100110011010000110010000100010001001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100100010001000110011001100110011001100110011001100110011010000110011001101000100010101010101010101010101010101010101010101100101010101010110011101110101010101110111011101110111011101110110011001100100010001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100111001110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110,
	2400'b001100110010001000100010001000100010001000100010001000100011001101000011010000110011001100110011001100100010000100010001000100100010001000110011001100110010000100010001000100010010001000100010001000100010001000100010001000110011001100110010001000110011001100110010001000100011001100110011001100110011001000100010001000100011001100110011001100110011010000110011010001000011010001000100010001010110010101010101010101010101010101100110010101010101011001110110010101100111011101110111011101110111011001110110010001000101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100111001110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011101110111011011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001100110100010001010101010000100010000100010001000100010010001000100011001100110011001000010001000100010001001000100010001000100010001100110010001100100010001000100010001100110010001000100010001100110011001100110011001100110010001000100011001100110011001100110011001101000100010001000100010001000011001101000100010101010101011101100110011001010101010101110110011001010101010101110110011001100111011101110111011101110111011101110111011001010100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100111011110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000010010010001000100010001000100001100100011001000100001000100010010001000100010001000110011001000010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000110010001000100011001100110011001000100010001100110011001100110011001100110011001100110011010001000100010001000100001100110101010001010101010101110111011001100110010101100111011001100110010101100111011001110110011101110111011101110111011101110111011101100101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100111011110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111011001100110011001100111011101100110011101110111011101110111011101110111011101110111011101110111,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000110100010000110011010000110010001000100001000100010001000100010001001000100010001000010001000100010001000100100010001000100010001000100010001100100010001000100010001000110011001100100010001000100010001100110010001000100010001000100011001000110011001100110011001100110011010001000100010000110100010001000100010101010101010101100111011101100110011001100111011101110110011001100111011101110111011101110111011101110111011101110111011101110111010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100111001110111011101110111011101110111011101110110111011101110111011101110111011101110111011101110111011101110111011011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110110011001100110011001100110011101110111011101110111011101110111011101110111011101110110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010000100010010010001000100001100110010001000100010000100010001000100010001001000010001001000100001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100011001100110011001101000100010001000100010001000100010001000100010101010101010101010110011101110110011101100111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100111001110111011101110111011101110111011101110111011011101110111011101110111011101110111011101110111011101110111011011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101011001100110011001110111011001100110011101100110011101110111011101110110011101110111011101100110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000010010000100010001001000110011001100110010001000100010000100010001000100010001001000100001000100100010001000010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000110011001100110011001100110100010001000100010001000100010001010101010101100101010101100101011001110110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110111110111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111011010100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100010001010101011001100110011001100111011101110110011101110111011101100110011101110111011101100110011001110110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010010001000100010001000100010001000010001000100010001000100010001000100010010001000100001000100010001000100010001001000100010001000100010001000100010001000100001000100100010001000100010000100100010001000100010001100110010001000100011001100110011001100110011010001000100010001010101010001000101010101010110010101100110011001110111011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110111101111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110111001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011001110110010001000100011001100110011001100110011001100110011101110110011001100110011001100111011001100110011001110110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000100001001000100010001000100010000100010001001000100010001000100010000100010001000100010001000100010001000100010001000100100010000100010001000100010001001000100010001000100001000100100010001000100010001000100001001000100010001000100010001000100010001000100011001000110011001100110011001100110100010001000100010001010101010101010101010101100110011001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101100111011101110111011101110111011101110111011011101111011011101110111011101110111011101110111011101110110111001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100110011101110111011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100100001101000101010101010101011001100110011001100110011001100110011001100110011101110111011101100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100001000100100010001000100010001000010001000100100001001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001000110011001100110100010001000100010001010101010101010110010101100110011001100110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011011111011101110111011101110111011101110111011101101110111011101110111011101110111011101110111011101110110101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011001110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101011001000011010001000101010101010110011001100110011001100110011001100110011001100111011101110110011001100110011101110110011001100110,
	2400'b001100110011001000100010001000100010001000100001000100100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110100010001000100010001000101011001010101011001100111011101100111011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011010110111101110111011101110111011101110111011101110111011101110110111011101110111011101110111101101110010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110110011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000100010000110100010101000101010101100101010101100110011001100110011001100110011001100110011001110110011001100110011101100110011001100110,
	2400'b010001000011001100110010001000100010001000010010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100011001000110011001100110011001000100010001000100010001000100011001100110010001100110011001101000100010000110100010101010100011001100101010101100111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001101111011110111011101110111011101110111011101110111011101110111011101110111011101101111011011101101010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110110010000110011001101000101010101000100010101010101011001100110011001100110011001100110011001100110011101100110011001110110011001100110011001100110,
	2400'b010101000100010000110011001100110011001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100001000100010001000100010001000100010001000100100010001000100010001000100010001000100011001100100010001000100010001000100010001000100011001100110011001100110011001100110100010001000100010001010101010101100110010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110111110111011101110111011101110111011101110111011101110111011101110111011011110111011011100100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100110011001101000101010001010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b010101010101010101000100010001000010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010101010101010001000110010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011100111011101110111011101110111011101110111011101110111011101110111011101110111011001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100111011101110111011101110111011101110110011101110110011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001101000101010001010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b010101100101010101010101010101000010001100100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100010010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001100100011001100110011001100110011001100110011010001010101010101000101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001110011101110111011101110111011101110111011101110111011101110111011101110110010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011001110111011101100111011101110111011101100111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110011001101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001100110011001100110010100110011010000110011001100100010001000100010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100001001000100010000100100010001000100010001000100010001000100010001000100001000100100010001000100010001000110010001101000011010001000011001100110011010001010110010101010101011001110110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100111001110111011101110111011101110111011101110111011101110111011101100101010011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101110111011101110111011001110111011101100111011101100111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110011001100110011010001010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001100110011101100110010001000101001100110100001100100010001000100010001000100010001000100010000100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100001101000100010101000011001101000110011001100110010101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011011110111101110111011101110111011101110111011101110110110111001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101100111011101110111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010001000011001100110011010001010101010001000100010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b010101100110011001100101010001010100001101000100010000110011001100100011001000100010001000100010000100010010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100100001000100010010001000100010001100110011001100100010001000100010001000100010001000100011001100100100001100100011010000110100011001010011010001000101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001101010111101111011101110111011101110111011011011101010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010001000011001100110011001101010101010001000101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001100110011001100100010001010100010001010100010001010100001100110011001000100010001000100010001000100010001000100001000100010001000100010001000100010001001000100001000100010001000100100001000100010001001000100001000100100010000100100010001000100011001100100010001000100010001000100010001000100010001100110011010001000010001101000100010101100100010001000100011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001101010111100110011001011101010101001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010000110011001100110011001101000101010001000100010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001010101010101010100010001010100010101010100010001000011001101000011001000100010001000100010001000100010001000100010000100010001001000100010000100010001000100100001000100010001000100010001000100010001000100100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100001101000100010001010101010001010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010000110011001100110011010001000101010001000100010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b011001010101010101010101010101000100010101000100010001000100001100110010001000100010001000100010001000100010001000100010001000010001000100100010000100010001000100010001001000100001000100010001001000010001000100100001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100011001100110100010001000101010001000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101100110011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010110011001110111011101110111011101110111011101110111011101110111011101110111011001100110010101010100010001000011001100110011010001010101010001000100010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b010101010101011001100110010101010101010101010100010001000100001100110011001000100011001000100010001000100010001000100010001000100001000100010001000100010001000100010001001000110001000100010001000100010010001000010010000100100010001000100010001000010001000100100001000100100010001000100010001000100010001000100010001000100010001000100011001100110100010001000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010110010101010111011101110111011101110111011101110111011101110111011101110110011001100110010101010100010000110011001100110011010001000101010001000101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b001100110011010001000101010101010100010101010101010101010100010001000100001100110011001000100010001000100010001000100010001000100010000100010001000100010001000100010001001001000011001000010001001000010010000100010010000100100010001000100010001000010001000100100001000100010010001000100010001000100010001000100010001000100010001000100010001100110011001101000100010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100101010101100101011001110111011101110111011101110111011101110111011101110110011001100110010101010100010000110011001100110011010001000100010001010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b001000100010001000100010001100110010001100110011010001000101010101010101010101000011001100100010001000110011001000100010001000100010000100010001000100010001000100010001000100110100001100100001000100010010000100010001000100010001001000100001001000010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001000100010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100111011001100101010101010110011001110111011101110111011101110111011101110111011101110110011001100101010101010100010001000011001100110011010001000100010001000101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000110011010001010101010101000011010000110010001100110011001100100010001000100010001000100001000100100010001000100010000100100100010000110001000100100010001000100001000100010001000100010001001000100001000100010001000100010010001000010010001000100010001000100010001000100010001000100010001100110011010000110011001100110100010001000100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101100111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100101010101010101011001100110011101110111011101110111011101110111011101100110011001010101010101010100010000110011001100110011010001000100010001000101010101010101010101010101011001100110011001100110011001100110011001100101011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000010010001000110100010001000100010001000011001100110100010000110010001000100010001000100010000100010010001100110011001000010011010100110001001000110010001100100001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001100110011001100110011001100110011001101000100010001000100001101000100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101100110011001100110011001010100010101010110011101110111011101110111011101110111011001100110011001010101010101000100010000110011001100110011010101000100010001000101010101010101010101010101011001100110011001100110011001010101010101010110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000010010001000100010001000100010001000100010001000100011010001000100010001000100001100100010001100100010001000100011001000100010001101000100001100100010010000100001001101000011010000100010001000100001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100111011101110111011101110111011101110110011101110111011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010110011001100110010101010101010001010110011001110111011101110111011101100110011001100110010101010101010001000100010001000011001100110100010101000100010001000100010001010101010101010101011001100110011001100110010101010101011001100110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000010010001000100010000100010001001000010001000100010010001000100011010001000100001100100010010000110010001100110100001100110010001001010100001100100001001000010001010001000011001100010010001000010001000100010001000100010001000100010001001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110110011101110111011001110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110010101010101010101010101010001000110011001100111011101110111011101110110011001100101010101010100010001000100010001000011001100110100010101000100010001000100010101000101010101010101011001100110011001100101010101010101011001100110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000100001000100010001000100010010001000010010001000110100001100100010001101000100010001000101010101000011000100110101010000100001000100010001001100110011001000100010001000010001000100010001000100010010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110100010001000100010001000011010001000100010001000100010001000101010001000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101000101011001010101010100110100011001100111011001110110011001100110010101010101010101010100010001000100010000110011001100110100010101000100010001000101010101010101010101010110011001100110011001010101010101010101011001100110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010000100100001000100010001000100010001000100010010001000100010001000100011010001000100010001000101010101010100001000100100010000100001000100010001001100100001001000100001000100010001000100010001001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000101011001100101010101000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001100111011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101010100010101100101010101000011010101010110011101100110011001100110010101010100010001000100010001000100010000110011001100110100010101000100010001000101010101010101010101100110011001100110010101010101010101010101010101010110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100001001000010001000100100010001000100010001000100010001101000100001100110100010101010101010000010011010100110001000100010001001000100010001000010001000100010001000100010010001000100001001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110100010001000100010001010101010101010100010001000100010001000100010001000100010001100111011101100101010001000101011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001100110011001100110011001100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100101010001000101010001000011010001000110011101100110011001100110010101010101010001000100010001000100001100110011001100110100010101000100010001000100010101010101010101100110011001100101010101000101010101000101010101010110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000010001000100100010001000100010001100100010001000100011001101010011001101010110010000100001010001000001000100010001001000010011001000010001000100010001000100010001000100010010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110100010001000100010101010101010101010101010001010100010001000100010001000100010001000101011001110111011001010100010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100110011001010101010101000100010001000100001101010101011001100110011001100110010101010101010001000100010000110011001100110011001100110100010101000100010001000101010101010101010101010110011001010101010001000101010001000100010001010110011001100110011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110010001001000101010100110101010101000001001101000010000100010010001000100011001000010001001000010001000100010010001000110011001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110100010001000101010101010101010101010101010101000101010101010100010001000100010001000100010101010110011101110110010101000101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110110011001110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001010101010101010100010001000100001101000101010101100110011001100110010101010101010001000100010000110011001100110011001100110100010101000100010001010101010101010101010101010101011001000100010001000100010001000100010101010101011001100110011001100110011001100101,
	2400'b001000100010001000100010001000100010001100100011001100100010001000100010001000100010001000100010001000100010001000110011010001010011001000100011010001010011010000110010001000110010000100010010001000110011001000010010001000010010001000100011010101000010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010101010101010101010101010101000101010101010101010101000100010001000100010001010101011001110111011001100101010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110110011001100110011001010101010101010101010000110011001100110100010101100110011001100110011001010101010101010100001100110011001100110011001100110100010101000100010001000101010101010101010101010101010101000100010001000100010001000100010001010101011001100110011001100110011001010101,
	2400'b001000100011001100110010001000100011001101000100001100100011001100100011001100110011001000100011010101000011010001000100010001000101010000100010001000110100001100110010000100100010000100010001000100110011000100010001000100010010001100110010001100100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001010101010101010101010101010101010101010100010001000101010101010101010101100111011101110110010101010100010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101100110011001100101010101010100010001000011001100110011010001010110011001100110010101010101010001000100010000110011001100110011001100110100010001000100010001000101010101010101010101010101010001010100010001000100010001000100010101010110011001100110011001100110011001010101,
	2400'b001100110011001100110011001000110011010101010101001100110100001100110011001100110011001100100100010101010100010101100101011001010100010101010100001000100010001000100010000100100001000100010001001000110010000100010001000100100010001000100010001100110100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001010101010101010101010101010101011001100111011001010110011101110111011101100101010001000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011001100110011101100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110110011001100110011001100101010101010100010001000100001100110011010001010110011001100101010001000100010001000100010000110011001100110011001100110100010001000100010001000101010101010101010101010100010001000100010001000100010001000101010101100110011001100110011001100110010101010110,
	2400'b001100110100010101000011001100110100011001100100001101000100001101000100001100110011001000100100010101010110010101100110011001110110010101010101010000100010000100010001000100010001000100010001001000100001000100010001000100010010001101000100010001010101010001000100010001000011001100110011001100110100001100110011010000110011001100110011010001000011001100110011001100110011001100110011001100110011001100110100010001010101010101100101010101100110011001010101011101110111011101110110011001010100010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100001110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101110111011101110110011001100110011001100101010101010101010101000100001100110011001101000101011001100110010101000100010001000100010001000011001100110011001100110100010001000100010001000100010101010101010001000100010001000011001101000100010001010101011001100110011001100110011001100101010101100110,
	2400'b001101010110010100110011001100110101011001010011010001010011010001000100001101000010001000100101010101010110011001100110011001110111011001100111011001010011000100010001000100010001000100010001000100010001000100010001000100010100011001100101010001000100010101010100010001000011001100110011010001010101001100110011010001010100001101000100010001000011010001000011001101000011001100110011001100110011001100110011001100110100010101010101010101010101010101000100011001110111011101110111011101100110010101000101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001111000100001111000100010001000100010001000100001110111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010001000100010001000101010101000100010001010101010101100110011001100110011001110111011001100110010101010101010101010101010001000011001100110011001100110100011001010101010101010100010000110011001101000100001100110011001100110100010001000100010001000100010001000100010001000100001100110100010001000101010101100110011001100110011001100110011001010101011001100110,
	2400'b010101110111010001000101010001010110011101010100011001010100010001000100010000110010000100110101010001100110011001100110011001100111011101100110011001000010000100010001000100010001000100010001000100010001000100010001000100010011010101100110010101000100010101000100010000110011001100110011010001000100001101000011010001010100001101000100010101000100010101000011010001000100010000110011001100110011001100110011001100110011010001000101010101010101010101010101010101100110011001110111011001100110011001010100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011001100111011001100110011001100110011101100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101111000011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101000100010001000011001100110011001100110011001100110011001100110011010001000101010101100110011001100110011001100110010101000101010101010101010101000100001100110010001000100100011001010100010101010100010000110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001010101010101100110011001100110011001100110010101010110011001100110,
	2400'b011001110110010001100101010001100111011101010110011001010101010000110100001100100010000100110100010101100110010101010101010101010100010000110010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001101000100001100110011001000100010001100110010001100110011010001000100010001000011010001010101001101010100010101010100010101010100010001010100010001000100001100110011001100110011001100110011001100110100010001010101010101010101010101010110011101110111011001110110011001100110010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010100010001000100010101010100010001000100001100110011001100110011001100110011001100110100010001000101011001100110011001100110010101010101010001000101010001000100010000110010001000100011010101010101010001000101001100110011001100110011001100110011001100110100010000110011001101000100010001000100010001000100010001000100010101010101010101010110011001100110011001100110010101100110011001100110,
	2400'b011101110100010101010101010101110111011001100110011001010100001100110011001000100001000100100011001000100010001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000110011001101000011010001100101001101010101010101100100010101010100010101010100010001000100010001000100001100110011001100110011001100110011010001000100010101010101010101010110011101110111011101110111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110110011101110111011101110111011001110111011101100110011001100111011001100111011101110111011101100110011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010001000100010001000101010101000100010001000011001100110011001100110011001100110011001100110011001100110011010001010110011001100110010101010101010001000100010001000100010000110010001000100011010001010100010000110100010001000011001100110011001100110011001101000101001100110011001101000011010000110100010001000100010001000100010001000101010101100110011001100110011001100101011001100110011001100110,
	2400'b011001010110011001010101011001110110011001110110010101000011001100100010001000100001000100010001000100010001000100010001000100010001001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010000100010001000100100010001000100010001000100010001000100010001000100010001000110011001100110100010001010101010101100101010101010100010101010100010001000100010001000100010001000011001100110011001100110011001101000100010001010101010101100110011001110110011001110111011101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100111011101110111011101110111011101110111011001110110011001100110011101110110011001110111011001100111011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101000101010101010101010001000100010001000100001100110011001100110011001100110011001100110011001100110011001100110011010001100110011001010101010001000100010001000100010001000011001000100010001101010100001100110011001101000100001100110011001100110011001101000100010000110011001100110011001101000100010001000100010001000100010001010101010101100110011001100110011001010110011001100110011001100110,
	2400'b010101100110010101100110011001110110010101010100001100100010000100010001000100010001000100010001000100010001001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110100010101100101010101010101011001010101010101000101010001000100010001000100010001000011001100110011001100110100010001000101011001010110011001100110011001110111011001100110011001100111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110110011001100111011101110110011001100111011001110111011101110111011101100110011001100110011001100110011001110110010101110111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101100110010101100101010101010101010101000100010001000011001100110011001000100010001100110011001100110011001100110011001100110011001100110100011001100110010101000100010001000100010001000011001100100010001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001010101010101100110011001100110010101010110011001100110011001100110,
	2400'b011001100101011101110110010101010100001100110010001000100001000100010001000100010001000100010001000100010010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010101010101011001100101011001010101010101000100010001000100010001000100010001000011001100110100010001000100010101100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011001100110011001100111011101100110011001100110011101110110011001110111011001100110011001100111011101100101010101110110011001100110011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110101011001100110011001010101010101010100010001000100010000110011010001000011001100110011001000100011001100110011001100110011001100100011001101010110011001010100010001000100010001000100001100100010001001000011001100110011001000110011001100110011001100110011001100110011001100110011001100110011010000110011010001000100010001000100010101010101011001100110011001100101010101100110011001100110011001100110,
	2400'b011001010110011101010101001100110010001000100010000100010001000100010001000100010001000100010001000100010001001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110100010101100101011001100101011001010100010001000101010001010101010101000100010000110100001101000100010001010110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011001100110011001110111011101100111011001100110011101110110011001100110011101100110011001110111011001110110011101100110011101110110011001010101010101100110011001100110011101110111011101110111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010110011001100111011001010101010101010101010101010101010001000100010001010101010001000100010000110011001100110010001000100010001000100010001000100100010101010101010001000100010001000100001100100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010101010101010101100110011001100101011001100110011001100110011001100111,
	2400'b011001010100001100100010001000100010001000010001000100010001000100010001000100010001000100010001000100010010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011010001000101011001100110011001100101010101000101010101010101010101010100010101000011001101000100010001000101011001100111011101100110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101100110011001110110011001100110011001100110011001100110011001100111011101110111011101100110011101100110010101010101010101100110011001100110011001110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110110011101110111011001110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001110111011001100110011001010110011001100100010001010101010101010101010101010101010001000011001100110010001000100010001000100010001000100010001101010101010001000100010000110011001100110010001000110011001100110011001100110010001100110011001100110011001000110011001100110011001100110011001100110011001100110011010001000100010101010101010101100110010101000101011001100110011001100111011101100110,
	2400'b010000110010001000100010001000100001000100010001001000010001000100010010001000100010001000100001000100100010001000100010000100100001001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001100100010001000100010001000100010001000100010001000110011001100110010001000100010001000100010001000100010001000100011001100110100010001010101011001100101010101010101011001010101010101100101011001010100010000110011001100110100011001100110011101100110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011001110111011001100111011001100110011001100110010101010110011101110111011101100111011101100101010101010101010101010110011001100110011101111000011101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110111011001100111011101100110011001100110011001100110010101010101010001000100001100110010001000100010001000100010001000100010001000100100010101000100010000110011001100110010001000110011001100100011001100100011001000100011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010101010101010101100101010001010110011001100110011101110110010101010110,
	2400'b001000100010001000100010001000100001000100010001001000100001000100010010001000100010001000100001000100100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001100110011001100100011001000100010001000100010001000110011001100110011001100100010001000100010001000100010001000100011001100110011010001000100010001010101011001100101011001100110011001100101011001100101010001000100001100110011010001100110011101100110011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110010101010110011001110111011101100111011101100101010101010101010101010110011001100110011101110111011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101100110011001100110011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110110011001100110011001010101010101010100010001000100001100110011001100100010001000100010001000100010001000100010001101000100010001000100001100110010001000100011001000100011001000100010001000100011001000100010001100110011001100110011001100110011001100110011001100110011010001000101010101010101010101010100010001100110011001110111011001000100011001100110,
	2400'b001000100010001000100010001000100010000100010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100100010001000010010001000100010010001000100010001000011001100110011001000100010001100110100010001000100001100110011001100100010001100110010001000100010001100110011001101000100010001000101010101010110011001100110011001100110011001110110010101000100010000110011001101010111011101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001010110011001100111011101110111011101100110010101010101010101010101011001100111011101110110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101100110011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100010001000100010001000011001100110011001000100011001000100010001000100010001000100010001000100011010001000100001100100010001000100011001100100010001000110011001000100010001000100010001000110011001100110011001100110011001100110011001100110011010001000101010101010101010101010100010101100110011101100100001101000110011001100110,
	2400'b001000100010001000100010001000100010001000010010001000010010001000100010001000100010000100100010001000100011001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000010001000100100010001000110100010001010101010001000101001100110011001101000100010001000100010000110011001100110011001000110011001100110011001100110011001101000100010001000100010101010101010101100110011001100110011001110110011001010100010001000011001101000110011101100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001010101010101100110011101110111011101100101010101010101010101100110011001100111011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100101010101010110011101100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010101010001000100010001000100001100110011001100110011001100100010001000100010001000100010001000100010001101000011001100110010001000100011001100100010001000100010001100100010001000100010001100110011001100110010001100110011001100110011001100110011010001000100010101010101010101000101011001100111010100110011010101100110011001100101,
	2400'b001000100010001000100010000100010010001000100010000100010010001000100010001000100010001000100010001100110011001100100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010000100010010001000100011010001010110011001000101011001000100010001000100010101010101010001000011001100110011001100100011001100110011001100110011001101000100010001000100010101010101010101010101011001100111011001110110011001100100010001010100010000110100011001100110011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010101011001100110011001100110011101100101010101100110011001110111011101110110010101010101010101010110011001110111011001010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110110011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101100110011001100110010101010100010001000101011001110110011101110111011101110111011101110111011101110111011101110111011001100110011001010110011001010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010101010101010100010001000100001100110100010000110011001100110011001000100010001000100010001000100010001000100011001100110010001000100010001000100010001000100010001000100010001000100010001101000011001100100011001100110011001100110011001100110100010001000101010101010101010001000101011001100100001101000110011001100110011001010100,
	2400'b001000100010001000100001000100100010001000100010001000100010001000100010001000100010001000100011001100110011001000100010001000010001000100010010000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001001000110011001100100010001010100010001000100010101010101010101000011001100110100010000110011001100110011001100110011001101000100010001000100010001000101010101010101011001100111011001100111011001100101010001010100010000110011010001100111011001110111011101100111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100101010101100101010101010101011001100110010101010101011001100111011101110101010101010101010101010101011001110110010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110111011001110111011101110111011001100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100101010101000100010001000100010001010110011001100110011001110111011101110111011101110111011101110110010101010110010101010110010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101010101010001000100010001000100010000110011001100100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000110011001000100011001100110011001100110011001100110100010001000101010101000100010001010110010100110011010101100110011001100101010001000100,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100011001100110011001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000010010001100110100010101100110001100110101010101010101010101010101010101010100010000110100010100110011001100110011001100110011001100110011010001000100010001010101010001010101011001100110011001100111011001100110010001000100010001000100001101000110011001100110011101100110011001100110011001100111011101110111011101110110011001100111011101110110011101110111011101100110011001100110011001100101010101010101010101010101010101010110011001010101010101100111011101100101010101010101010001010101010101010101010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011001100110011101100110011001110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011001100101010001000100010000110011010001000101011001010110011101100110011001100110011001100111011101100110010101010101010001010101010101010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110010101010101010101010101010000110100010101000100010000110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001100110011001100110011001100110100010001000100010001000100010101100101001101000101011001100101010101010101010001000011,
	2400'b001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110010001000100010001000100001000100100001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001100110011001101000101010101000100010101010101010101010101010101010100010101000100010101000011001100110011001100110100001100110011010001000100010001010101010101010101010101010110011001110110011001100110010101010100010001000100001100110100011001100110011001100110011001100110011101100110011101110111011101110110011001100110011101110111011101100110011001100110011001100110011001100110011001100101010101010110010101010101010101010110010101010110011001100110010101010101010101010110010101010101010101010101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110110011001010101010101010100001100110011001101000100011001010101011001100101011001100110011101100110010101010101010001010100010001010101010101010101011001110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101010101010101010100010001010100010001000100010000110011001100100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001100110011001100110011001100110011010001000100001100110101011001000011010101100110011001100101010001010100010001000011,
	2400'b001000100010001000100010001100100010001000110010001000100011001100110011001100110100001100100011001100100010001000100001000100100001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100100010001100100010001000100010001000100100010000110011010001000100010001000101010001010101011001010101010101010100011001010011001100110011001100110011001100110100010001000100010001000101010101010101010101010101011001110110011001100110011001010100010001000100010101000011010001100110011001100110011001100110011001100110011001110110011001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010001000101010101010110011001100110010101010101010101010101010101100110010101010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101100110011001100111011101110111011001100111011101110111011101110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101000100010000110011001100110100010101010100010101100101011001100110011101100101010001000100010001000100010101000100010101010110011001110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101010101010101000100010101010101010101010100010000110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100011001100110011010000110100010001000011010001010110001100110101011001100110010101000100001101000100001100110011,
	2400'b001000100010001000100010001100100010001000110011001100110011010001000100001100110100001100110011001000100010000100010001000100010001001000010001000100010001000100010001000100010001000100010001000100010001000100100011010001000011001100110010001000100010001000100011010001000100001100110011010001000100010101010101011001010101010101010101011001100100001101000011001100110011001100110011010001000100010001000100010101010101010101010101010101100111011001100110011001010101010001010100010001000011001101010110011001100110011001100110011001100110011001100110011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010001000100010101100101010101100110010101000100010101000100010101010101010101010101011001100110010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011001110111011101100111011001110111011101110111011001110111011101110111011101110110011101100111011101110111011101110111011101110111011101110110011001110110011001100110010101000100010001000011001100110011010001000011010001010101010101100110011001100101010001000100010001000100010001000100010101100111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101100110010101010101010101010101010101010100010001000011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001100110011001000100010001100110010001100110011010001000100001100110100010101100100010001010110010101100100001100110011001100110011001100110011,
	2400'b001000100010001000100010001100110011001000110011001100110100010001000100010001000100001100110011001000100010001000010001000100010010001000010001000100010001000100010001000100010001000100010001000100010001000100100011010001010100001101000011001000100010001000100010001101000100010001000011001100110011010001010101011001100101011001100101011001100101001101000100010000110100001100110011001101000100010001000101010101010101010101010101010101100110011001100110011001100101010101010101010101000100001101000101011001100110011001100110011001100110011101100110011001100111011101110111011001100110011001100110011001100110011001100110011001110110011001100110011001100110010101010101010001000100010001010101010101010101010101000100010001000100010001010101010101010101010101010101010101100110011001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011101110111011101110111011101100111011101110111011101110111011101110111011001100111011101110110011101110111011101110111011101110110011001110110011001100101010101000100010001000100001100110011001101000011001101000100010101010110011001100101010001000100001101000100010001000101010101100110011101110111011101110111011101110111011101100111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001010101010101010101010101010101010101000011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000011001001000101010101010101011001100101010101000011001100110011001100110011001100110011,
	2400'b001000100010001000100010001100110011001000110100010000110100010001010101010101000100001100100010001000100010000100010001000100010010000100010001000100010001000100010001000100010001000100010010000100010001000100100011010001010110010001000100010000100010001000100010001001000100010001000100010000110011001101000101010101010101011001100101011001100101010001000100010000110011001100110011001100110011010001000101010101010101010101010101011001100110011001100111011101100110011001010110011001010100010001000100011001100110011001100110011001100110011001100110011001110111011101110111011101110110011001100110011001100110011001100110011001100111011001100110011001100110011001010101010101000100010001000100010101000100010001000100010001000100010001010101010101010101010101010101011001010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001110110011001100110011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101100111011001100110011001100110010101010011010001000100001100110011001100110011001100110100010001010101011001010100010001000011001101000100010001000101010101010110011101110111011101110111011101110111011001110110010101100111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100101011001010101010101100110010101000100010000110011001100110010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001100110010001000100010001000110010001000100011001100110010001101010101010101010101011001010100001100110011001100110011001100110011001100110011,
	2400'b001000100011001100110010001101000100001100110100010000110101010101010110010101000100001100100010001000100010000100010001000100100010000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001010110011001000100010100110010001000100010001000110100010101010101010000110011001100110011010001010110011001100110011001100110010001010100010000110011001101000011001100110011001101000100010101010101010101010110011001100110011001100110011101100110011001100110011001100101010001010100010001100110011001100110011001100110011001100110011001100110011001100110011101110111011001100110011001100110011001110111011001100110011001100111011001100110011001100110011001000100010001000100010101010100010001000100010001000100010001000101010101010101010101010110010101010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101100110011001110111011101100111011101110111011101100111011101100110011101110111011101110111011101110110011001100110011001100110010101010100001100110011010000110011001100110011001100110011010001000101010101010100010001000011001101000100010001000101011001100110011001110111011101100111011101100110011001010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101100110011001010101010101100101010101010101010001000011001100110011001100100010001000100010001000100010001000100010001000100001001000100010001000100010001000100010001000100010001101000011001000100010001000100010001000100011001100100011010101010101010101010101010000110010001000110011001100110011001100110011001100110011,
	2400'b001100110011010001000010010001010100001100110100010001000101011001010110010101000100001100100010001000100010000100100001000100100010000100010001000100010001000100010001000100010001000100010001000100010001000100100011010001010110011001100100010001000011001000100010001000100011010001010110010100110011010000110011001101000101011001100110011001110110010101010101010001000100001101000011001100110011001100110100010001010101010101010110011001100110011001100110011001100110011001100110011001100110010001100101010101010110011001100110011001100110011001100110011001100110011001100111011101110111011101100110011001100110011101110111011001100110011001100110011001100110011001100110011001100100010001000100010001010101010001000100010001000100010101010101010101010101010101010110010101010110010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101100110011001110110011001100110010101100101010000110011001100110011001100110011001100110011001101000100010101010100010000110011001100110100010001000101010101100110011101100110011101110111011001010101010101010101011001100110011001110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011001100110011001010101010101010101010101010011001101000100001100100010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000100010001000110010001000100010001000100010001000100011001000110100010101010100010001000011001000100010001000100010001000100011001100110010001100110011,
	2400'b001100110100010001000011010001010101010001000100010101000101011001100101010001010100001000100010001000010010001000100001001000100001001000010001000100010001000100010001000100010001000100010001000100010001000100100011010001010101011001100110010001000011001000100010001000100010001101010101010101010011010001000011001100110100010101100110011001110111010101100101010101010100010001000011001100110011001100110011010001010101010101010110011001100110011001100110011001100110011101110110011101100110010101010110011001000101011001100110011001100110011001100110011001100110011101100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110010101010110011001100110010001000100010001000101010101000100010001000101010101010101010001000101010101010101011001010110011001010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101011001110111011101110111011101110111011101110111011101110110011001110110011001100110011001100110010101000011001100110011001100110010001000110011001100110011010001010100001100110011001100110100010001000101010101010110011001100110011001100110010101010101010101010101010101010110011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001010101010101100101011001000100010101010100001100110011001000100010001000100010001000100010001000100010001000100010001000010001000100100010001000100010001000100010001000100010001000100010001000110011001101000100010000110011001000100010001000100010001000100010001000100011001100110011001100110011,
	2400'b010001000100010101010101010001100110010001000101011001010110011001010100010101010011001000100010000100010001000100010001001000010001001000100001000100010001000100010001000100010001000100010001000100010001000100100011010001000101011001100111011001000011001100100010001000100010001001000101010101010101010001000101010000110011010001010110011001110110010101100101010101010101010001000100001100110011001100110011001101000101010001010110011001100110011001100110011001100110011101100110011001100110011001100110011001100100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001010101010101010110010101000100010001000100010101000100010001000100010001000100010001000101010101010101010101100101010101010110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101000100010001000100010001010101011001110111011101110111011101100110011101110111011001100110011001100110011001100101010101010100001100110011001100100010001000100011001100110011001101010100001100110100010000110100010001000101010101010110011001100110011001100101010101010101010101010101010101100110011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101100110010101010101010101010100010001000011001000100011001000100010001000100010001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001100100011010001000011001100100010001000100010001000100010001000100010001000100010001100110011001100110011,
	2400'b010001000100010101010101010101110111010001000110011001010110010101010110010101000011001000100010001000100010001000100010000100010001000100100001000100100010000100010001000100010010001000010001000100010001000100100011010001010101010101100111011101100100001100110010001000100010001000100100010101010101010000110100010101000011001101000110011001110110011001100101010101010101010001000100001100110011001100110011001100110100010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110010101000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010100010001000101010101010101010001000100010001000100010001000100010001010100010001000100010101010101010101100110010101010110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100101010101000100010001000100010001000011010001000101010101100111011101110110011101110111011101110111011001100110011001100110011001100110011001010101010000110011001100110010001000100011001100110011001101000011001100110100010001000100010001000100010101010101010101100110011001010101010101010100010001010101010101100110011101110111011101110110011001100110011001100101010101010100010001000100010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100101010101100110010101000100010101000011001100110011001000100010001000100010001000100010001000010010001000100010001000100010001000100010001000100010001000100010001000100011001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011,
	2400'b010001000101010101010110011001110111010101000111011101100101010101100101010101000011001000100010001000100010001000100010000100010001001000100010000100010001001000010001000100010010001000010001000100010001000100100011010001010101011001110111011101110110001100100010001000100010001000100011010001010101010101000011010101010100001101000100010101010110011101110110010101100101010101010100010000110011001100110011001100110100010101100110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001010101010101010101011001100110011001100110011001100110011001100110011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010101010101010101010101010001000100010001000101011001110111011101110111011101110111011101100110011001100110011001010101010101010101010001000011001100110011001000100011001100110011010000110011001100110011001101000100010001000100010101010101010101010101010101010100010101000100010001010101010101100110011101110111011001100110011001100101010101000100010001000100010001010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011101100101011001100110010101010101010000110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011,
	2400'b010101010101010101100110011001111000011001010111011101010110011001100101010100110011001000100001000100010001001000100010000100100010001000100010001000010001001000010001000100010001001000100001000100010001000100100100010001010101011001110111011101110110010000100010001000100010001000100010001101000110010101010011010001010100010000110011010001000101011001110111011001100101010101010100010001000011001100110011001100110011010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001010101010101010101011001100110011001100111011001110111011001110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011001100101010101000100010001000100010001000100010001010110011101110111011101110111011101110110011001100110011001100110010101010101010001000011001100110011001100100011001100110011001100110011001100110011001101000100001100110100010101010101010101010101010101000101010001000100010001000100011001100110011101110110011001100110010101000100010001000100010001000100010001000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110110010101010101010101000100010001000100001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001000100010001000100010001100110010001000100011001100110011,
	2400'b010101010101011001100110011101111000011001010111011001010110010101010101010000110010001000100001001000100001001000010001001000100010001000100010001000010001000100010001000100010010001000100001000100010001000100100100010101010101011001100110011001100101010000110010001000100010001000100010001000110101010101100101010001010101010101000011001101000101010101100111011001100110010101100101010001000011001100110011001100110011010001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110010101100101010101010101010101010101010101010100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001010101010001000100010001000100010001000100010001100111011101110111011101110111011001010110011001010101010101010100001101000011001100100011001100110010001100100011001100110011001100110011001100110011001100110100010001010101010101010100010101010100010001000100010001010101011001100110011001100110011001010100010001000100010001000100010001000101010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011001110110010101010100010001000100010001000100001100110011001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001101000100,
	2400'b010101100110011001100111011101111000011001100111011101010110010101010100010000100001000100100010001000010010000100010010001000100001001000100010001000100001000100010010001000100001000100100010001000010001000100100100010101010110011001100111011001100101010101000011001000100010001000100010001000100011010101100110010001000101010101000100010001000100010001010111011101110110010101010101010001000100001100110011001100110011010001000100011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110011001100110011001100110011001100101010101010101010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010110011101110110011001110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101010101010101000100010001000101010001000101011001110111011101110111011101100110011001100101010101010100001100110011001000100010001100110010001100100011001100100011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010101010101011001100110011001100101010001000011010001000100010001000101010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011001100110011001100101010101010100010000110011001100110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110100,
	2400'b010101100110011101110111011110001000011001101000011001010110010101000011001000010010001000100010001000010010001000010010001000100010001000100010001000100010001000100010001000100010000100010001001000010010000100110101010101010110011001100111011001100101010101000100001000100010001000100010001000100010001101010110010101000101010101010100010001000100010001010110011101110111011001100101010101000100001100110011001100110100001101000100010101100110011001100110011001110110011001100110011001100110011001100110011001100110011001100111010101100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110011001100110011001100110011001100101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100110011001100110011001010101010101000100010001000100010001010101010101010110011101110111011101100110010101010101011001010101010000110011001000100010001000100010001000100011001100100011001000110011001100110011001100110100010001000100010001000100010001000100010001010101010101000100010101100110010101000011001100110011010001000101010101010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010101010001000011001100110100001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010001000100001100110010001000110010001000100010001000100010001000100010001000110010001100110011001100110011010001000100,
	2400'b011001110111011110000111100010001000010101100111011001010100010000110010000100100010001000010010001000100010001000100010001000100010001000100010001000100010001000010010001000100010001000010001000100010010001000110101011001100110011001100111011001100101010101000100001100100010001000100010001000100010001000110101011001000101010101010101010001000100010001010101011001110111011001100110011001010101001100110011001100110100001101000100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101100110011001100110011001100101011001010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001100110011001010101010101010101010101000100010001000101010101000101011001110111011001100111011001010101010101000100001100110011001100100010001000100010001000100010001100110010001000110011001100110011001100110100010001000100001101000100010001000100010101010101010101010101011001100100001100110011001100110011010001000100010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010100010001000100010001010100001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001000101010101010101010000110010001000100010001000100010001000100010001000110011001100110011001100110011001100110011010001000100,
	2400'b011001110111100010000111100010001000010101110111011001000100010000110001000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000010001001000100001001000100010001000100010001101000101011001100110011001110111011001100101011001010101001100110010001000100010001000100010001000100011010101100100010101000101010101000100010001000101010101100111011101100110011001100110010001000011001100110011001101000100010001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101010101010101010100010001000100010001000100010001100111011001100110011001100101010001000011001100110011001000100010001000100010001000100010001000110010001100110011001100110011001100110100010001000011001101000100010001000101010001010101010101100110010101000011001100110011001100110011010001000100010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100111011001100110010101010101010101000100010001000100010000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101010110011001010100001100100010001000100010001000100010001000100010001100110011010001000100010001000100010001000100010001000100,
	2400'b011001110111100010000111100010000111010101110111010101000011001100100001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000100100010001000100010001000100011010101100110011001100111011101110111011001010110010101010110001101000010001000100010001000100010001000100010010001100101010101100101011001010100010001000101010101010111011101110110011101110110010001000100010000110011010001000100010101010110011001100110011001100110011001100110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110010101100101010001000100010101010100010001000100010001000100010001000100010001000101010001010100010001000100010001010101010101100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001010110010101010101010101000100010001000100010101000110011101100110011001100110010101000011001100110010001000100010001000100010001000100010001000100011001100100011001100110011001100110100010000110011001101000100010001000100010001010110011001010100001100110011001100110011001100110011001100110100010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110111011001100110011001010101010101010101010101000100010001000100010001000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001100110010101000011001000100010001000100010001000100010001000100011001100110100010001000100010001000100010001000100010001000100,
	2400'b011101111000100010001000100010000110010101110110010001000011001000100010001000100010001000010001001000100010001000100010001000100010001100100010001000100010001000100010000100010010001000100010001000100100011001100111011001110111011101110110011001100101010101100110010001000010001000100010001000100010001000100010001000110101011001100101011001100101010001000101010101010110011101110111011101110110010101010100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110010101010100010001010101010101010101010101000100010001000100010001000100010001000101010101010101010001000101010101010101010101010110011001100110011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100101010101010101010001000100010001010101010101100110011001100110011001010100001100100010001000100010001000100010001000100010001000100011001100110011001000100011001100110011001100110011001101000100010001000101011001100110010101000011001100110010001000100011001100110011010001000101010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101010101010101010101010100010001010100010001000011001000100010001000100010001000100010001000100010000100010010001000100010001000100100010101100101010000100010001000100010001000100010001000100010001000100011001101000100010001010101010001010101010001010101010001000100,
	2400'b011110001000100010001000100010000101011001110101010000110010001000100010001000100010001000010010001000100010001000100010001000100011001100100010001000100010000100100010001000100010001000100010001000110110011101110111011101110111011101110111011001100110011001110110010100110011001100110010001000100010001000100010001000100011010101100110010101100101010101000100010001010101011001110111011101110111011001010101010101000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011101100110011001100110011001100110011001100110011001100110011001100110010101010100010101010101010101100101010101000100010001000100010001000100010001000100010101010101010101000100010101010100010001010110011001100111011101110111011001100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010101010101010101010101000100010001000100010001010110011001100110011001010101010000110011001000100010001000100010001000100010001000100010001101000011001100100011001100110011001100110100001101000100010001000101011001010101010000110011001100110011001100110011001101000100010101010101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101010101010101100110010101010101010101010100010001000100010001000011001000100010001000100010001000100010001000100010000100100010001000100010001000110101011001010101001100100010001000100010001000100010001000100010001000110011010001000101011001010101010101000101010101010101010101010100,
	2400'b011110001000100010001000100010000101011101110101001100100010001000100010000100100010001000100010001000100010001000100010001000100011001100110010001000100010000100010010001000100010001000100010001001000110011101110111011101110111011101110111011001100110011001110110010000110100010001000011001000100010001000100010001000100010001101010110010101100110010101010101010101010101011001100111011101110111011101100110010101010100010001000100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110011001100101010001000101010101010101011001010101010001010100010001000100010001000100010001000100010001010101010101010101010001010101010101010110011001100111011001110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101010110011001010101010101010101010101000100001101000101011001100110011001010101010100110010001000100010001000100010001000100010001000100010001100110011001100110010001100110011001100110100001101000100010001010101010101000011001100110011001100110011001100110011001101000100010101010110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100101010101010101010101010101010101010101010101000100010001000100010000110011001100110011001000110010001000100010001000100010001000100010000100010010001001010110011001010011001000100010001000100010001000100010001000100010001100110100010001000100010101010100010001010100010001010101010001010101,
	2400'b011110001000100010001000100001110101011101100011001000100010001000100001000100100010001000100010001000100010001000100011001100110011001100110010001000100010001000100010001000100010001000100010001101010111011101110111011101110111011101110111011101100111011101110110010000110100010101010100001000100010001000100010001000100010001000110110011001010110011001010101010101010101010101100111011101110111011101100110011001010100010001000100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100110011001100110011001100110011001100110011001100110011001100101010101010101010101010110010101010101010101000100010001000100010000110100010001000100010001000101010101010101010101010101010101010101011001100111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101111000100001110111011110000111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010110011001100110010101010110011001010101010101010100010000110100010101010110010101010110010101000011001000100010001000100010001100110011001100110011001100110011001100110010001100110011001100110011001101000100010101010101010100110011001100110011001100110011001100110100010001000100010001010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001010101010101010101010101010100010101010101010101000100010001000100001100110100010000110011001100110010001000100011001100110010000100100010001000010001001001000101010001000011001000100010001000100010001000100010001000100011010001010100001100110011001101000100010001000100010001000101010101010101,
	2400'b100010001000100010001000100001010110011001000010001000100010001000100001000100100010001000100010001000100010001000100011001101000100001100110010001000100010001000100010001000100010001000100010001101100111011101110111011101110111011101110111011101110111011101110110010001000101010101010101001100100010001000100010001000100010001000100100011001100101011101100101010101010101010101100111011101110111011101100110011001100101010001000100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101100110011001100110011001100110011001100101011001100110010101010101010101010101010001000100010001000100001100110011010001000100010001000100010101100110010101010101010101010101011001100111011001110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101100111011101100101011001100110011001100110011001100101010101000011010001000110010101000100010001000100001100100011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001101000100010001000101010000110011001100110011001100110011001101000100010001010101010101010101011001010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110010101010101010101010101010101000100010001000100010001000100001100110100010001000100010001000011001101000100010001000011000100100010001100100010001001000011010001000010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011010001000100010001000100,
	2400'b100010001000100010001000011101010110010100110010001000100010001000100010001000010010001000100010001000100010001000110011010001000101010000110011001000100001000100100010001000100010001000100011010101110111011101110111011101110111011101110111011101110111011101110110010101010110011001100101001100100010001000100010001000100010001000100011010001110110011001100101010101010101010101010110011101110111011101100110011101100101010001010100010001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101100110011001100110011001100110011001100110011001100101010101010101010101000100010001000100010001000100010000110011010001000100010001000100010001010110011001010110011001010101011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001110111011101111000100010001000100010000111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101100111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101100110011101100110011001010101010101010100010001000100010101010011010001010100001100100010001000100010001100110010001000110010001000100010001100110010001100110011001100110011010000110100010001000011001100110011001100110011001100110011001100110011001101000100010001010101010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010101010101010100010001000100001100110100010001000100010000110011001101000100010000110011001100110011001100110011001000100001001100110010001000100011010000110010001000100010001000100010001000100011001100100010001000100010001100110011001100110011001100110011001100110011001100110011,
	2400'b100010001000100010001000011001010101010000100010001000100010001000100010001000100010001000100010001000110010001100110011010001000101010000110011001000100001000100100010001000100010001000100100011001110111011101110111011101110111011101110111011101111000011101110110011001100110011001100110001100110010001000100010001000100010001000100010001101010111011001100110010101100101010101010101011101110111011101110111011101100110010101010101010001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011001100110011001100110011101100110011001100110011001100110011001100101010101000101010001000100010101000100010001000100010001000011010001000100010001000100010001000101011001100110011001100101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011110000111011110001000011101110111011101111000100001110111011110001000100010001000100010001000100001111000011110001000100001111000100010001000011110000111011101111000100001110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101100110011001100110011001010101010101010101010000110011001101010100001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000110011001100110100010001000011001100110011001100110011001100110011001100110011001101000100010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100101010101010101010101010100010001000100010001000100010001000100010001000011001100110011001000100010001000010010001000100010001000010001001000110010001000100011001100100010001000100010001000100010001000100010001000100011001100100011001100110011001100110011001100110011001100110011001100110011,
	2400'b100010001000100010000111010101010100001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001000101010000110100001000100010000100100010001000100010001000110110011101110111011101110111011110001000011101110111100010000111011101110111011101110111011101110110010000110010001000100010001000100010001000100010001000110110011001100110010101010110010101010110011001110111011101110111011101110110010101010101010001000101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011001100110011001100110011001100110011001100110011001100110011001010101010001000100010001000101010101000100010001000100010001000100010001000100010001000100010001000101010101100110011101100101011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000011101111000100010000111011101111000100001110111011101110111011101111000100001110111100001110111011101111000100010001000011110000111011110000111011101110111100001110111011110001000011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110110011001100110010101010101010001000100010000110011001100110100010000110010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001101000100010000110011001000110011001100110010001100110011001101000100010001000100010101010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001010101010101000100010101010101010001000100010101010100010001000100010001000011010001000011001100100010000100010001000100010001000100010001000100100010001000100011001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011010001000100010001000100010001000100,
	2400'b100010001000100001110101010001000011001000100010001000100010001000100010001000100010001100100010001000110011001100110011010001000101010000110100001000100010001000100010001000100010001001000111011101110111100010001000100010001000100010001000100001110111100010000111011101110111011101110110010001000011001000100010001000100010001000100010001100110100011001100110011001100101011001100110011101110111011001100111011001110111011001100110010101000100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110110011001100111011101100110011001110111011101110110011001100110011001100110011001100110010101010100010001000100010001010101010001000100010001000100010001000100010001000100010001000100010001000100010101010110011001100110011001100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010001000100010000111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010000111100010001000011110001000100010001000011110001000100001110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111011101100111011101100110010101010101010101000100010000110011001100110011010001000011001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011010001000100001100100011001100110011001100110011001100110011001100110011010001000100010001010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100101010101010101010101000100010101000100010101010100010001000100010001000100001100110011001000100010001000010001000100010001000100010001000100010001001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110100010001000100010101010101010101010100,
	2400'b011101110110011001010101001100100010001000100010001000100010001000100010001000100011001100100010001100110011001100110011010001010101010101000101001100100010001000100010001000100010001001000111011101110111100010001000100010001000100010001000100001111000100010001000011110001000100001110110010101000011001000100010001000100010001000100010001000100011010001100110011001100110011001100110011001100111011101100111011101110111011001100110010101000100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110110011001100110011001110110011001100110011001110111011001100110011001100110011001100101010101010100010001010100010101100101010001000100010001000100010001000100010001000100010001000100010001000100010001010110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101110110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010101000100010001000100001100110011001101000011001000100010001000100010001000100010001000100010001000100010001000100010001000110010001100110011010001000011001000100011001100110011001100110010001100110011001100110011010001000100010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001010101010101010101010001000100010000110011001100110011001000100010001000100001000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001100110011001100110011001100110011001100110011001100110011010001000100010001000101010101010101,
	2400'b011001010110011001100100001000100010001000100010000100100010001000100010001000100011001100110010001100110011001100110011010001010101010101010101001100010010001000100010001000100010001001010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001010011001000100010001000100010001000100010001000100010001101000101010101100110011001100110011001100111011101110111011101110111011101100110011001010100010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100111011101100110011001100110011001110110011101100110011001100110011001100110011001100110011001100101010101010100010101010101011001100101010001000100010001000100010001000100010001000100010001000100010001000100010101010101011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100001111000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010101010101010101010001000100010001000011010000110011001100110010001000100010001000100010001000100010001000100010001000100011001100110010001100110011001100110011001000110011001100100010001100100010001000110011001101000100010001010101010101010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110010101010100001100110011001100110010001100110010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010010001000100011001100110011001100110011001100110011001100110011001101000100010001010101010101010101010101010101,
	2400'b010101010101011001010011001000100010001000100010001000100010001000100010001000110011001100110010001101000100001100110011001101010101010101010100001000010001000100100010001000100010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100100001100110010001000100010001000100010001000100010001101000100010101100110011001100110011001100110011101110111011101110111011101100110011001100100010001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011001100110011001110110011101110110011001100110011001100110011001100110011001010100010001000100010101010110011001010100010001000100010001000100010001000100010001000100010001010101010101010100010101010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011001100111011001110110011101100101010101010110011001010100010001000100010001000011001100100010001000110011001000100010001000100010001000100010001000100010001000100010001100110010001000110011001100100011001000100010001000100010001000100010001101000100010001000100010101010101010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110010101000011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010010001000010001000100010001000100100010001000100010001000110011001100110011001100110011001100110100010001000100010001000101010101010101010101010101,
	2400'b011001010110010100110010001000100010001000100010001000100010001000100010001000110100001100110011001101000100001101000100001101010101011001010101001100100010001000100010001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110101001100110010001000100010001000100010001000100010001100110100010101100110011001100110011001100110011101110111011101110111011101100110011101100101010001010111011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101110111011001110111011101100110011001100110011101110111011001100110011001100111011001100110011001000100010101000101011001100110011001010100010001000100010001000100010001000100010001000100010001010101010101010101010101010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011001100110011101100110011101110111011101110111011001110111011101110111011101110111011101110111011001100110011001100110011001100110011001100111011001100111011101110111011001110111010101110111011001010101010101100110011001010100010001000100010000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110010001000100010001000100010001100110011010001000100010101010101010101010101011001100110011001100110011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110110011001000011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001100110011010001000100010001000100010101010101010101010101010101010101,
	2400'b011001100101010000100010001000100010001000100010001000100010001000100010001000110100001100110011001101010101010001000100010001000101011001100100001000100010001000100001001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101110101001101000011001000100010001000100010001000100010001000110011010001010110011001100110011001100110011001110110011001110111011101110110011101100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110110011001100111011101100110011101100111011101100110011001100111011001100110010001000101010001010110011001100110011001000100010001000100010001000101010001000100010001000100010001000101010101010101011001010101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010000111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110110011001110111011101110111011101110111011101110110011001100110011101100110010101010101010101010101010101010101010101100101011001100110011001010101010000110100010001000100010001010101010101000100010000110011001100110010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000110010001000100010001000100010001000100011001100110100010001000101010101010101010101100110011001100110011001100111011001100110011001100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001010100001100100010001000100010001100110011001000100010001000100010001000100010001000100010001000010010000100010001000100010001000100010001000100010001000100010001000100010001000100100010001000100010001000100010001000100010001000100010001000110011001101000100010001000100010101010101010101010101010101010101,
	2400'b011001010101001100100010001000100010001000010010001000100010001000100010001001000100010001000011010001010101010001000101010001000101011001100100001000100010001000100010000100100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110101010001010011001000100010001000100010001000100010001000100011010001010110011001100110011001100110011001110111011101110111011101110110011101110110011001010110011001100110011001100110011001100110011001100110011001100110011101100111011001110111011001110111011101110111011101110111011101100111011101110110011001110111011001100110011001100110011001100101010101010100010101100110011001100110010101010100010001010100010001010101010001000100010001000100010001000101010101100101011001100101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010000111011110001000011110001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011001100111011001110110011001100111011101110111011101110111011101110111011101110111011001110111011101100111011101110111011101110110011001100110011001010101010101010101010001000101010001000100010001000100010101000100010001000011001100100010001000110100010101010101010000110011001100110011001000100010001000100010001000100010001000100011001000100010001000100010001100110010001000100010001000100010001000100010001000110011010001000100010001000101010101010110010101100110011001100111011001010101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100101010000110010001000100010001000110011001100110010001000100010001000100010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001100110100010001010101010101010101010101010101011001100101,
	2400'b011001010100001000100010001000100010001000100010001000100011001000100010001101000101010001000100010001010110010101000101010101000101011001010011001000100010001000100010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101110101011001100100001000100010001000100010001000100010001000100010001101000101011001100110011001100110011001110111011101110111011101110110011101110110011001010110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011001100110011101010101010101010101010101100110011101110110010101010101010101010101010001010101010001000100010101000100010001000101010101100101010101100110010101010110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010101011001010101010101010101010001000101010001010100010001000100001100110011001100110011001000100010001000110100010000110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001000100011001100110100010001000100010001010101011001100110011001010110011001100101010101010101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110010101000011001000100011001100110011001100110011001000100010001000100010001000100010001000100010001000100011001100100010000100010001000100010001000100010001000100010001000100100001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000110100010001010101010101010101010101010101011001100110,
	2400'b010101000010001000100010001000100010001000100010001000100011001000100011001101000101010001000100010001010110011001000101010101000101011001010011001000100010000100010010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100001100111100010001000100001100101011101110100001000100010001000100010001000100011001000100010001100110101011001100110011001100110011001110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100111011001100110011001100111011001010101010101010101010101100111011101110101010101010101010101010101010001000100010001000100010101000100010001000100010101010101010101100111010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110011001100110011001100101010101010100010101010101010101010101010101010100001101000100010000110011001100100010001000100011001101000011001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100010001100110011001100110100010001010101011001100101010101010101010001000100010001000100010001000101010101010101010101100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101001100100010001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100011001100110010000100010001000100010001000100010001000100010001000100100010000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000110011010001010101010101010101011001100110011001100110,
	2400'b010100110010001000100010001000100010001000100010001000110010001000100011001101010110010101000100010001100110011001010101011001010100011001010011001000100010001000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000011101100110011101110101001100100010001000100010001000100011001100100010001000110100011001110111011001100110011001100111011101110111011101110111011101110110011001100101011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011001110111011001110110010101010101010101010110011001100111011101100101010101010101011001100101010001000100010001000101011001010100010001000100010101100101010101100111011001010101011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110110011001100110011001100110011001100110010101010101010101010101011001010110011001100100010101100101010001000100010000110011001000100010001000100011010001000011001100110100001100110010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000110011001101000101011001010110011001010100001100110011001100110011001100110011010000110011010001000100010101010101010101010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001100110011001100110011001100110011001000100010001000100011001100110011001100110010001000100010001000100010001000010001000100010001000100010001000100010001000100010001000100010001000100010001001000100001001000100010001000010010001000100010001000100010001000100010001101000101011001100110011001100110011001100110,
	2400'b001100100010001000100010001000100010001000100010001100110010001100110100010001010110010101000101010001100111011101010101011001100100011001010011001000100010001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100111011101110101001100110010001000100010001000100010001100110010001000110011010101100111011101100110011001100111011101110111011101110111011101110111011001100101011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100111011101110110011101100101010101010101010101010110011001100111011001010110010101010101011001100101010001000100010001000101011001010100010101000101010101100110010101100110011101100101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011101110111011101100101010101010101010101010110011101100111011101010101010101010100010001000100010001000100001100110010001000100010001101000100010001000100010001000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110100010101010110010101000011001100100010001000110010001000100010001100110011001100110011001100110100010001000101010101010101010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010000110010001000100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010010000100100010001000100010001000100010001000100010001000100010001000100010001000110100010101100110011001100110011001100110,
	2400'b001100100010001000100010001000100010001000100010001100110011010000110101010001010110011001010101010101100111011101100101011001100110010101010011001000100010001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001111000100001110100010001000011001000100010001000100010001000110010001000110011010001100110011101110111011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101100110011001010101010101010101011001100110011101100111011001100110010101010110011001110101010101010100010001010110011001100101010101010101010101100110010101100110011101100101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010110011001010110011001100111011101100110010101010101010001000100010101010100010001000100010001000011001100100010001000100011010101010101010101010101010000100010001000110011001000100010001000100010001000100010001100100010001000100011010001000100010001000011001100100010001000100010001000100010001000100011001100110011001100110011001100110011010001000100010001010101010101100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100100001100110011001100110011001100110011001100110011001100110011001100110100001101000100010101010100010000110011001100110010001000100010001000100010001000010001001000100010001000100010001000100010000100100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101010101011001100110011001100110,
	2400'b001000100010001000100010001000100010001000100011001100110011010101000101010001010110011001010101010101100111011101110101011001100111010101010011001000100010001000100010001101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001111000100001110100010101000011001000100010001000100011001000110011001000100011010001010110011101110110011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001010101011001010110011101100111011101110111011001100110010101010110011001110110010101010101010001010111011101100101010101010101011001100110011001100110011101110110010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110110011001100110011001100110011001100110011001100110011001100110010101100110011001010101010101000100010001000100010000110011001000100010001101010110010101010110010101000010001001010101001100110010001000100010001000100010001100100010001000110011010001000011001100100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110100010001010101010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001100110011001100110011001100110011001100110011010001000100010101010101010101010101001100110011001100110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000010010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010101100110011001100110,
	2400'b001000100010001000100010001000100010001000100011001100110100010101000101010001010111011001100101010101100111011101110110011001100111011001000011001000100010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011110001000100001100101011001010100001100100010001000100011001100110011001100100011001101000110011101110111011001100111011101110111011101110111011101110111011001100110011001100110011001100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101100110011001100110011101100110011101110111011101110110010101100110011101110110010101010101010101100111011101100101010101010101011001100111011001100110011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101011001110110011001100110011001100110011001100101010101010100010101010101010101010100010001000100010001000100010001010100010000100010001000100100011001100111011101100100000100110110001101000100001100110010001000100010001000100011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100011001000110011001100110011001100110011001101000100010101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010100110011010000110011001100110011001100110011001100110011001100110100010001000101011001010101011001100101010000100011001100100010001100110011001100100010001000100001001000100010001000100010001000100010000100010010001000100011010000110010001100110010001000100010001000100010001000100010001000100010001000100010001000100011001101010101011001100110,
	2400'b001000100010001000100010001000100010001000110100001100110101010101000101010001000111011101100101010101100111011101110111011001110111011101000010001000100010001000100011010110001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100001110111100010001000100001100110011001100101001100100010001000100011001100110011001100100010001100110101011001110111011101100111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011001110111011101100110011101110111011101110110010101100110011101110110010101010101011001110111011101110110011001010110011001100111011001100110011001110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110110011101100110011001010101010001000100001100110011001101000011001100110011001101000100010001000100010001000100010001000100001100100010001101100110011001100110001000100101001101010101010101010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101001100110100001100110011001100110010001100110011001100110100010001000101010001010110010101100110011001100101010100110010001000100010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100011010001000011001101000011001100110011001000100010001000100010001000100010001000100010001000100010001000100011010101100110,
	2400'b001000100010001000100010001000100010001101000100001100110101011001010101010001000111011101110110011001100111011101110111011101110111011101010011001000100010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000011101100111011101100110010000100010001000110011001100110011001100110010001100110100011001110111011101100111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100111011101110111011101100111011101110111011101110110010101100110011101110111010101010110011101110111011101110110011001010110011001110111011101100111011001110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110110011001100101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000010000100100101011001100110001100010100001001000101010100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010000110011001101000101010101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001000011010001000100001100110011001100110011001100110011001101000100010101000110011001010110011001100101010101010101010001000011001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001000100010001000100010000110010001000100011001000100010001000100010001000100010001000100010001000100010001101010110,
	2400'b001000100010001000100010001000100011001101000100001101000101010101010110010001000110011101110110011001100111011101110111011101110111011101100011001000100010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000011101100111011101110111010000100010001000100011001100110011001100110011001100110100010101100111011101100111011101110111011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011001100111011101110110010101010111011101110111011101110110011001100110011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010001000100010001000100010001000100010001000100010001000100010101000101010101010101010101010101010101000101010001000011010001000100001100100010010001100101001100010010001000110100001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011010001000100010000110100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111010100110100010001000100001100110011001100110011001100110011001101000101011001100110011001100110011001100110011001010100001000100010001000100010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100011010001000100010001000100001100100010001000110011001000100010001000100010001000100010001000100010001000100010001000110100,
	2400'b001000100010001000100010001000100011010001000100001101000110010101010110010101000110011101110111011001110111011110000111011101110111011101100011001000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001110111011101110111010000110010001000100010001100110011001000110011001100110100010001010111011101100111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011001100111011101110110010101100111011101110111011101110110011001100110011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010100010001000100010001000100010001000100010101000100010001000101011001010110011001100110011001100101011001100110011001010101010001000011001100110001000100110100001100100001000100100010001000100010001000100010000100010010001000100010001000100010001000100010001000110010001100100010001100110011010001000100010001000100010001000100001100110011001100110011001101000100010001000011001101000101011001110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101100101001101000100010001000011001100110011001100110100001100110100010001000110011001100110011001100110011101100110011001100101001100110010001000100010001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010101000100010101000011001000100010001100110010001100110010001000100010001000100010001000100010001000100010001000100011,
	2400'b001000100011001000100010001000110100010101000100001101000110010101010110011001000101011101110111011101110111100001110111011101111000011101110100001000010001001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100001110111010101000011001000100011001100110100001000100011010001000100010001000110011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101100110011101110110011001110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101010101010101010101010101011001010101010101010101011001100110011101100111011001100101011001100110011001010110011001100101010000110010000100010010001100100010001000100001001001010011001000100010001000010010001000100010001000010010001000100010001000100010001100110010001100110100010001000101010101010101010101000100010001000100010000110011001100110011010001000100010000110100011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011010001000100010000110011001100110011001100110100010001000100010001000100011101110111011101110110011001100110010101010101010000110011001000100010001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010101010101010000110010001000110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010,
	2400'b001100110011001100100010001000110101010101000100010001010110010101010110011001000101011101110111011101110111100010001000011101111000100001110101001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010000111010101010011001000110011001100110100001100110011001101000100010001000101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110110011101110111011001110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101100110011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101010101010101010101010110010101010110011001010110010101100110011001110111011001100101011001100110010101010100010001000100010001000101010101010100001000010010001000100001000100010010010101100100001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010101000101010101010101010101010100010101010100010001000011001100110011001100110100010001000100010001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111010101000100010001000100001100110011001100110011001101000100010001000100010001010100010101111000011101110111011101100101010101000100010000110011001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010101010100001100110011001101000011001100110100001100110010001000100010001000100010001000100010001000100010001000100010,
	2400'b001100110011001100100010001101000110010001000100010001010110010101010110011101010101011110000111011101111000100010001000100010001000100010000101001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001110111100010001000100010000111011001100100001100110011001100110100001100110011001101000100010101000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110011001100111011101100111011101110111011101110110011001110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101010101010101010101010101100110010101100110011001100110011001100110011001100111011101110111011001010100010001000011001100110011001100100010001000100010001101000100010000100001000100010001000100010100011001100011001000100010001000100010001000100010001000100010001000100010001000100010001101000011001100110100010101010110011001010101011001100101011001100101010101100101001101000101010000110011010001010100010001010110011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001110101010001000011010001000011001100110010001100110011010001000100010001000101010101100110011001100111011101110111011101100101010001000100010001000011001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000110101011001010101010101010101010101010100010001000011010000110011001100100010001000100010001000100010001000100010001000100010,
	2400'b001100110011001100100010001101010110010001000100010001010110010101100110100001100101011110001000100001111000100010001000100010001000100010000101001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010000111011101110101001100110011001100110100010000110011001100110100010101010100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001100111011001100111011001110111011001110111011101110111011101110111011101110110011101100111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101010101011001010110011001100110011001100110011001100110011001100110011101100110011001010101010000110011001100110010001000100010001000100010001000100010001000100010010001000011000100010001000100010010001100110010001000110010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010101100110011001100110011001100110010101100110011001100110010101010110011001100101010001010110011001010101011001110111011101110111011101110111011101110111011101110110011001100111011101110111011101100100001100110011010000110011001100110011001100110100010001000100010101010101010101100111011101100111011101110111011001100101010101010100010001000010001000110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100101011001100110011001010101010101010101010101000100010000110100001100110011001100100010001000100010001000100010001000100010,
	2400'b001100110011001100100010010001100110010001010100010101100110010101100111100001110101011010001000100010001000100010001000100010001000100001110100000100100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110101010000110011001100110100010100110011001100110100010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011001110111011001100110011001110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010000110011001100110011001100100010001000100010001000100010001000100010001000100001001000110100001000010001000100010001000100010011010000110011001100110011001100110011001100100010001000100010001000100010001000100010001100110100010001010101011001100110011001100110010101100110011001100110011001100110011001100110010101010110011101100101010101100111011101110111011001100111011101110111011101110111011001100110011101110111011001000011001100110011001100110011001100110011010000110100010101000101010101010110011001100111011101110111011101110110011001100101010101010101010001000010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011001100110011001100110011001100110011001010101010001000100010001000100001100110011001000100010001000100010001000100010,
	2400'b010001000011001100100011010101100101010001010100010101110110010101110111100010000110011010001000100010001000100010001000100010001000100001110100001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110101010000110011001100110100010100110011001100110100010101010101010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110011001110110011001100110011001100110011001100110011101110111011101110110011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101010101011001100110011001100110011001100110011001110110011001100110011001100110010101010101010001000100001100110011001100110010001000100010001000100010001000100010001000100010001000010001001000010010001000010001000100010010001000100100010001010100010001000011001100110011001100110011001100110011001000100010001000100010001000100011001100110100010101010110011001100110011001100110011001100110011001100110011001100111011001100110011101110110010101010110011101110111011101110111011101110111011101110111011101100111011101110110010000110011001100110011001100110011001100110100010001000100010101010101011001010110011101110111011101110111011101100110011001100101010101010101010000110010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100100011001100110011001100110011001100110011001010101010101010100010101010101010001000011001000100010001000100010001000100010,
	2400'b010001000011001100110011010101110101010101010101010101110101010101110111100010000111011001111000100010001000100010001000100010001000100001110011001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110010100110011001100110100010101000011001100110100010001010110010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100110011001100111011101100110011001100110011001100110011101110110011101110110011001110111011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100101010101010100010001000100010000110011001100110011001100110010001000100010001000100010001000100010001000100010001000100001000100010001000100010001000100010001000100100010001101000101010000110011001100110011001100110011001100110011001100110010001000100010001000100010001000110011001101000100010001010101011001100110011001100110011001100111011101110111011101110110011001110111011001100101011001110111011101110111011101110111011101110111011101110111011101110100001100110011001100110011001100110011001101000100010101000100010101010101011001100110011101110111011101110111011101100110011001010110011001100101010100110011010001000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110101011101110111011101110111011001100110011001100110011001010101010101100101010101000100001100100010001000100010001000100010,
	2400'b010001000011001100110100011001100100010101010101011001110101010101110111100010001000011001111000100010001000100010001000100010001000100001100010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100001110111011101110110010101000011001101000100010101000011001101000100010101010110010101010111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011101110110011001110111011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001010101010001000100010001000100010001000100001100110100001100110011001100100010001000100010001000100010001000100010001000100011001000100001001000010001000100010001000100010001001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100100010001000100010001000110011001100110011001100110100010001000101011001100110011001100110011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101010011001100110011001100110011001100110011010001010100010101010100010101010101011101100111011101110111011101110111011001100110011001100110011001100110010100110011010100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100101011001110111011101110111011101110110011001100110011001100101011001100110010101010101001100110011001100100010001000100010,
	2400'b010101000011001100110100011001100100010101010101011101110101010101110111100010001000011101111000100010001000100010001000100010001000100001010010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100001110111100001110111011001000011010001000101010101000011001101000100010101010110011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111100001110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110110011101110111011101110111011101110111011101110111100001110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110110011101110110011001110111011001110110011101100110011001110110011001110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100101010001000100010001000101010101000100010001000011001101000100001100110011001100100010001000100010001000100010001000100010001000100010001000010010000100010001000100010001000100010001000100010010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110100010101010110011001110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110110011101110111011000110011001100110011001100110011001100110100010001010101010101100101010101100110011101110111011101110111011101110110011001100110011001100110011001100101001100100011010000110100010000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011010101110111011101110111011101110110011001100111011001100110011101110110011001100101010000110011001100110010001000100010,
	2400'b010101000011001100110101011101100101011001010101011101110101011001110111100010001000100001111000100010001000100010001000100010001000100001000010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100001110111011001000100010001000101010101010011001101000110010101010101011001010101011101110111011101110111011101111000100010000111011101110111011110001000100010001000100010001000100010000111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110110011101110111011101110111011101110111100010001000100010001000100010001000100001110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011110000111100010001000100001111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110110011101100110011001110111011001110111011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011001100110011001100110010101000100010001000100010101010101010101010101010000110100001100110100001100110011001000100010001000100010001000110010001000100010001000100010000100010001000100010001000100010001000100010001000100010010001000100011010001010101010000110010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001101000011001101000100010101100111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110110010000110011001100110011001100110011001101000100010101010101011001010101011001110110011101110111011101110111011101110111011001100110011001110111011101110101001100110011010101010100001100110010001000100010001000100010001000100010001000100010001000100010001000110011001100110011010001010110011101110111011101110111011101110110011001100111011101110110011001100101010001000011001100110011001000100010,
	2400'b010000110011001101000101011101110101011001100110011101110101011110000111100010001000100010001000100010001000100010001000100010001000011100110001001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010000111011101010100010001000101010101010011001101000110011001100101010101010101011110001000100001111000100001110111100010001000011110001000011110001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100111011101110111011101111000011101110111100010001000100010001000100010001000100010000111100010000111011101110111100001110111100010000111011110000111100010000111100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011001100110011001110110011001100110011001100110011001110111011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110110011001010101010001000100010001000100010101010101010101010101001100110100001100110100010000110010001000100010001000100010001100110011001000100011001000100010000100100010001000010001000100010001000100010001001000100010001000110110011101110110011001010011001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001000011001100110011010001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100110011001100110011001100110011010001000101010101100101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110110001100100100011001010011001101000011001000100010001000100010001000100010001000100010001000100010001000110011001100110100010101010110011001110111011101110111011101100111011101110111011101110110011001100110010101000100010000110011001100100010,
	2400'b010000110011001101000101011101110110011101100110011110000110011110001000100010001000100010001000100010001000100010001000100010001000011000100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010101010101000101010101010011001100110101011001110111011001010101011010000111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101100110011101110111011101110101011101111000011101100111011101110111011110001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100001110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101100110011001100110011001100111011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101010001010101010101010110011001000011001100110011001101000100001100110010001000100010001000100011001100110011001100110011001100100010001000010001000100010001000100010001000100010001001000100010001000100101100001110111011101010011001100100011001100100011001000100010001000100010001000100010001000110011001101000011001100110011010001000011001100110011010001000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011010000110100001100110011001101000100010001010101011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100100101011001010011010000110010001000100010001000100010001000100010001000100010001000100010001100110011001100110100010101100110011101110111011101111000011101111000011101110111011101100110011001100110010101010100010001000100001100110010,
	2400'b010000110011010001000110011101110110011101110111011110000110011110001000100010001000100010001000100010001000100010001000100010001000010100100001001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100110010101010101010101010100001100110100011001110111011101100101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110110011001111000100001110110011010001000011101100111100010000111011101110111011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010000111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101100110011101100110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010101010101010101010001010101011001100110010100110011010000110011010001000011001100110011001100110010001100110011001101000100001100110100001100100010001000010001000100010001000100010001000100010001001000110011001100100010011010001000011101010100001100110011001100110011001100100010001000100010001000100010001000100010001000110011001101000100001100110011001100110011010001000100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110100001101000100001100110011010001000100010101010101011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001100110110011001000011001100100010001000100010001100110010001000100010001000100010001000100011001100110011001100110100010001010110011101110111011101111000100010001000100001110111011001100111011101110110011001010100010101000100010000110011,
	2400'b010001000100010001010110011101110111011101110111011110000111011110001000100010001000100010001000100010001000100010001000100010000111001100100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001010101010101010100001100110100011001111000100010000111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100111011110000110011010001000011001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001111000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100111011101110111011001100111011101100111011001100110011101110111011101110110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100101010101010110010101010100001100110011001100110011010000110011001100110011001100110011001100110011001101000101010000110011001000100010001000100001000100010001000100010001000100010001000100100011001100110011001101101000011101010100001101000011001101000011001100100010001100110010001000100010001000100010001000100010001100110100010001000011001100110011010001000100010001010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010000110100010001000100001100110011010001000100010101010110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110110010100110011001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000100010001010101011001110111011101111000100010001000100010000111011101110111011101110111011001010101010101010101010001000011,
	2400'b010001000100010001010110011101110111100010000111011110000111100010001000100010001000100010001000100010001000100010001000100010000111001000100001001000110111100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001010110010101010100001100110100011001111000100010000111011001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100110011110000110011010000111011001110111011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101100111011101110111011001110110011001100111011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010101011001010110010101000011001100110011001100110011001101000011001100110011001101000011001100110100001101000101010000110010001000100010001000100010001000010001000100010001000100010001000100100011001100110011001100110110011101010011010001000100010001000011001100110100001100110010001100110011001000100010001000100010001000100011010001000100010000110011010001000100010001000110011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100010001000011001100110100010001000101011001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001001000110010100110011001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000100010101100110011001110111011101111000100010001000100001110111011101110111011101110111011001010110010101010101010101000100,
	2400'b010001000100010001100110011110001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010000101001000010001000101001000100010001000100010001000100010001000100001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001010110011001010100001100110100010101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001100111011101110110010101110110011001110110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011001110111011001100111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110110011001100110010101000101010101010101010000110011001100110011010000110011001101000011001100110011001101000100001100110100010001000100001100110011001000100010001000100010001000010001000100010001000100010001000100010010001101000011001100110011011101100101010001000100010101010100001101000100010000110011010000110011001100100010001000100010001000100010001000110100010000110011010001000100010001000100010101110111011101110111011101110111011101110111011101110111011101110111011101110100010001000100010001000100010001000100010001010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001001000110010000110011001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110100010101100110011101110111100010001000100010001000011101110111100001110111011101110111011001110110010101100101010101000100,
	2400'b010101000100010101100111100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001001011000100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101100110011001010100010001000100010101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001100110011101100110010101100101011001100110011001100110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100001110111011101111000100010001000100010001000100010000111011101110111011101110111011101110110011101110110011001110111011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110010000110100010001000100001100110011001100110100010000110011001101000100010001000100010000110101010100110100001100110011001100110011001000100010001000100010001000010001000100010001000100010001000100010001001000110100010000110011001101100110010101100101010101010100010101010101010001000101010001000011001100110011001100100010001000100010001000100011010001010100001101000100010001000100010001010111100001110111011101110111011101110111011101110111011101110111011101010100010001000100010001000100010001000100010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001101000101001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000100010001010110011101110111100010001000100010001000100001110111011101110110011001110111011101110110011001100101010101000100,
	2400'b010101010101010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001001101000100010001000100010001000100010000111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101100111011001010100010001000100010101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100101011001100110010001010101011101100101010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100100001100110011001101000100001100110011001100110100001101000100010001000101010001010100010001000101010101000011001100110011001100110010001000100010001000100010000100010001000100010001000100010001000100010001000100100011010001000100001101000110011101110110011001100110011001100101010001010100010101000100010001000011001100110010001000100010001000100010001101000100010001000100010001000100010001000101011101110111011101110111011101110111011101110111011101110111011001000100010001000100010001000100010001000101010101100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001101000100001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000101010101100110011001110111011101111000100010001000100010000111011101110111011101110111011101110110011001100110010101000101,
	2400'b010101010101010101100111100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100001100010001000100001001001111000100010001000100010001000011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101110111011001010100010001000100010101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100101010101100101010001000110011001010110010101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001000011001100110011010001000011001100110011001101000011001101000101010001010100011001100101010001000100010000110011001100110011001100110010001000100010001000100001000100010001000100010001000100010001000100100001000100010010001101000100010000110011011001110110011101100110011001100101010101010101010101000100010001000100001100110011001000100010001000100010001000100011010101010100010001000100010001000100010101110111100010000111011110000111011101110111011101110111010001000100010001000100010001000100010001010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001101000100001100110010001000100010001000100010001000110010001000100010001000110011001100110011001100110100010001000100011001110111011101110111100010001000100010001000100010001000100001110111011101110111011101110110011101100110010101010101,
	2400'b011001100101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001101111000100010001000100010001000011101110111011110001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011001111000011001010101010001000100010101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100101011001010100010001000101010101010101011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110100010001000011001100110011010001000100010001000101010101010101010101100110011001100100010000110011001100110011001100100010001000100010001000100010000100100001000100010001000100010001000100010001000100010001001001000100010000110011010001100111011101100111011001100101010101010101010101010101010101000100001100110011001100110011001000100010001000100011001101010101010001000100010001000100010001100111011101110111011101110111011101110111011101110110010001000100010001000100010001000100010101100110011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011001101000011001100110010001000100010001000100010001100110010001000100010001000110011001100110011001100110100010001010101011001110111011110001000100010001000100010001000100010001000100001110111011101110111011101110110011101110110010101010110,
	2400'b011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010010110001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000011001010101010001000100010101101000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100101010001000100010001000101010101100111011101111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100001100110011001100110100010001000011001100110011010001000100010001000101010101100110011001100110011001100101001100110011001100110011001000100010001000100010001000100010001000100010000100010001000100010001000100010001000100100010001000100100010001000011001001010111011101110111011101100110011001010101010101010101010101000100010001000011001100110100001100100010001000100011001100110100010101000100010001000100010001000110011101110111100001110111011101110111011101110100010001000100010001000100010001000100010101100110011101110111011101110111011101111000011101110111011101110111011110000111011101110111011101110111011101110111011101110111011101100011001101000011001100110010001000100010001100110011001100110010001000100010001000110011001100110011010001000100010101010110011001111000100010001000100010001000100010001000100010001000100001110111011101110111011101100111011101110110010101100110,
	2400'b011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010011010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000011101010110010001000100010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110010101010110010000110100010001000100010101100111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000011001100110011001101000100010001000100001101000100010001000100010001010110011001100111011101110111011001010011001100110011001100110010001000100010001000100010001000100010001000100010000100100010001000010001000100010010001000100010001000100011010001000100001100110110011101110111011101110110011001100110011001010101010101010101010001000100010001000100001100110011001100100010001000110011010001010100010001010101010101000100010101111000011101110111011101110111011101100100010001000100010001000100010001010101011001100111011101110111011110000111100010001000100001110111011101110111100001110111011101110111011101110111011101110111011101110111011101100011010001000011001100100010001000100011001100110011001101000010001000100010001000110011001100110011010001000100010101100110011001110111011110001000100010001000100010001000100010001000011101110111011101110111011101110111011101110101011001100110,
	2400'b011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100110010101000101010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100110010101000101010000110011001101000100010001010101011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001000110011001101000100010001000100010001000100010001000100010101010110011001100111011101110111010101000011001100110011001000100010001000100010001000100010001000100010001000100010000100010001001000010001001000100010001000100010001000100010001101000100001100110100011101110111011101110111011001100110011001100110011001100101010101000100010001000011001101000011001100110010001100110011001101000100010001000101010101010101010101100111011101110111011101110111011101010100010001000100010001000100010101010110011001110111011101110111011110001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011010000110011001100100010001000110011001100110011010001000011001000100010001000110011001100110100010001000100010101100110011001110111011101111000100010001000100010001000100010001000100010001000100001110111011101110111011101100110011001100110,
	2400'b011101110110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111010000100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100111010101010110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110011001100101010001000100010000110011001100110100010001000110100001110111100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100011001100110011001100110011010001000100010001000100010001000100010101010101010101100110011101110110011101110110010000110011001100110011001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010000110011010101111000011101110111011101110111011001100110011001100110010101010100010001000100010001000011001100110011001100110011001100110100010001000101010101010101010101010110011101110111011101110111011101010100010101000100010001000101010101100110011101110111011101111000100010001000100010001000100010000111011101110111011101111000011101110111011101110111011101110111011101110111011101010011010000110011001100100010001000110011001101000100010001010011001000100010001000110011001100110100010001000100010001100111011001110111100010001000100010001000100010001000100010001000100010001000011101110111011101110111011001100110011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000110001100100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100101010101100101010001000100010000110011001100110100010001010110011101100111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001100110011001100110100010101000100010001000101010001010101010101100110011001100111011101110110011001010100001100110011001100110010001000100010001000100010001100110011001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100011010000110011010001101000100010000111011101110111011101110111011101110110011001100101010001000100010001000100001100110011001100110011001101000100010001000100010101010101010101010101011001110111011101110111011001000100010101010100010101010101011001100111011101110111011101111000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101010100010000100011001100100010001000100011001101000100010101100100001000100010001000110100001100110100010001010101010001100111011101110111100010001000100010001000100010001000100010001000100010000111011101110111100001110111011001110111011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110010101010100010001000100010001000100001101000100010001010111011001100111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110011001100110011001100110101010101000100010001000101010101010110011001100110011001110111011101110111011001010100010000110011001000100010001000100010001000100011001100110011001000100010000100100010001000100010001000100010001000100010001000100010001000100010001000100010010000110011001101011000100010000111011101110111011101110111011101110110011001100110010101000101010101000100010000110011001100110011001101000100010001000100010001010101010101010101010101100111011101110111010101000100010101010101011001100110011101110111011101110111011110001000100010001000100010000111100010000111100010001000011110000111100001110111011101110111011101110111011101110111011101000100001100100011001100100010001100110011010001000101010101010011001000100010001000110100010001000100010001010101010101010111100001110111100010001000100010001000100010001000100010001000100010001000100001111000011101110110011101110111011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111100010001000100001110111011101100110010101010100010001000100010001000011001101000100010001010110010101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010011001100110011001100110011001101000110010101010101010101010110010101100110011001100110011101110111011101100110010101000100010000110011001000100010001000100011001100110011010001000011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001101000111100010001000100010001000100001110111011101110110011001100110010101010101010101010100010000110011001100110011001101000100010001010101010101010100010101010101010101010110011101110111010101000101011001010110011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000011110000111011101110111011101110111011101110111011101110111011101000100001100100011001100110010001100110011010001000100010101000010001000100010001000110100010001000100010101010101010101010111100010000111011110001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110011001100110011001010101010101100111011101110111011001010101010001000100010001000100010001000011001100110100010001010101010101100110011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110011001100110011001100110011010001010110010101010101010101010110011001110111011101110111011101110111011101010101010101000101010000110010001000100010001100110011001100110100010101000100001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001101000110100010001000100010000111100001110111011101110110011101110111011001100110010101010101010101000011001100110011010001000100010001010101010101010101010101010101010101010110011101110110010001010110011001100111011101110111100001110111011101110111100010001000100010001000100010001000100010001000100010000111011110000111011101110111011101110111011101110111011101110111011001000011001000110011001100110011001100110100010001000101010101000010001000100010001000110100010001000100010101010101011001100111100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110000111011101110111011101110111,
	2400'b011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011001010101010101010101011101110110010101010101010001000100010001000100001100110011001101000100010001010101011001100111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001100110011001100110011010001000101010101100111011001100101011001100110011101110111011101110111011101110111011101100100010001010100001100100010001000100011001100110011001101000101010101010100001000100010001000100010001000100011001100100010001000100010001100110011001100100010001000100010001000100010001101000110011110001000100010001000100001110111011101100110011101110111011101100110011001100101010101010100001100110011010001010101010001010110010101010101010101010101010101100110011101110110010001100111011001110111011101110111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011101110111011101110111011101110111010101000011001000110011001100110011001100110100010101010101010101000011001000100010001000110100010001000101010101010101011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111,
	2400'b011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011001100101010101010101011001110110010101010101010001000100010001000011001100110011001101000100010001010101011001100111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101000011001100110011001100110100010001010110010101110111011001100110011001100111011101110111011101110111011101110111011101100100010001000011001100100010001000110011001100110011010001010110011001010011001100100010001000100010001000110011001100110011001000100011001100110011001100100010001100110011001100100010001001000101011110001000100010001000100001110111011101100111011101110111011101110111011001110110011001010100001100110011010001010101010101010101010101010101010101010101010101010110011001100101010001100111011101110111011101111000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111010101000011001000110011001100110011001100110100010101100101011001100101010000100010001000110100010101010101010101010110011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111,
	2400'b011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111011101100110011001100110010101100110011001100101010001000100010000110011001100110011001101000100010101010101011001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010000110011001100110011001101000101010001100110011001110111011001100110011101110111011101110111100010000111100001110111100001100011001100110011001000100010001000110011001100110100010101100110011001010011001000110011001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100100010001000110100011110001000100010001000100010000111011101100111011101110111011101110111011101110111011001100101010000110011010001000110011001010101010101100101010101010101010101010101010101010100011001100111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110110010001000010001100110011001100110011001101000100010101100110010101100110010100100010001000110100010101010101010101100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111,
	2400'b011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100110011001100110011001010110011001010100010001000100001100110011001100110011001101000100010101010110011001110110011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001101000011001100110100010001010110010101100110011001110111011101110111011101110111011110001000011110001000100001110111011101100011001100110011001000100010001000110011010000110101011001100111011001010011001000100010001000100010001000110100010001000100010001000011001101000011001100110011001100110011001100100010001000100100011110001000100010001000100010001000011101110111011101110111011101110111011101110111011101110110010100110100010001000110011001100101011001010110011001100101011001100110010101010101011101100111011101110111011110001000011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010000111011110001000100001111000011110000111011101110101010101000011001100110011001100110011001101000101011001110111010101010110001100100010001000110100010101010101011001100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110011001100101010101010100010001000100001100110011001100110011001101000100010101010110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000011101111000011101111000100001110111011101110111011101110111011101110111011101110111011101110111100001010011010001000011001101000100010001100110010101110111011110000111011101110111100010001000100010001000100001111000011110000111011101110100001100110010001000100010001100110011010001000101011001110111011001010011001000100010001000100010001100110100010001000101010101010100010001000100001100110011001100110011001100110010001000100011011001111000100010001000100010001000100001110111100010000111100001110111011101110111011101110111011001000100010001000101011001110110011001100110011001100110010101100110010101010110011101110111011101110111011101111000011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100100010100110011001100110011001100110100010001000101011001110111011101100110010100100010001000100100010101010110011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010000100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100111011001100101010001010100010001000100001100110011001100110011001101000100010101100110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101111000011101000100010001000100010001000100010101110110011001110111011110000111011101110111100010001000100010001000100010001000100010000111011101110100001100110011001000100011001100110011010001010110011001110111011001010011001000100010001000100010001101000101010101010101011001010100010001000100001101000100001100110011001100110011001000100010011010001000100010001000100010001000100010001000100010001000100001111000011110000111011110000111011101010100010101000101011001110111011001010110011001010110011001100110010101010110011101110111011101110111011101110111011101110111100010001000011101111000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000011101100101010100110011001100110011001101000100010001000101011101110111011101110111010100100010001000100011010101100110011001100110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100101010001000100010001000011001100110011001100110011001101000100010101010101011001100110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101111000011110000111010101000101010101000100010101010101011001110110011101110111100010001000100010001000100010001000100010001000100010001000100010000111011101110100001100110011001100110011001100110100010001100111011101110111011101010100001000100010001000100010001101010101011001100110011001100100010101010101010001000100010001000011001100110011001000100010010110001000100010001000100010001000100010001000100010001000100010001000011110000111100010000111011101110110011001000100010101110111011101100110011001100110011001100111011001010110011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000011101010101010000110011001100110100001101000100010101010110011101110111011101110111010100100010001000100011010101100110011001100110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101010100010001000100010001000100001100110011001100110011001101000101010001000100010001010101010101100111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010101010101010101010101010101010101011101110110011110000111100010001000100010001000100010001000100010001000100010001000100010000111011101100011001100110011001100110011001100110100010101110111011101110111011101100100001000100010001000100011010001010110011001110111011001100101011001100110010101010100010001000100001100110011001000100010010001111000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100001110111011101010101010101100111011101100110011001100110011001100111011001100111011101110111011101110111011101110111011101110111011101111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010101010000110011001101000100010001000101010101100111011101110111011110000111010100100010001000100011010101100110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100000100100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001010100010001000100010001000100001100110011001100110011001100110011001101000100010001000100010101100110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101010101010110010101100101010101010101011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101000011001100110011001100110011001101000100011001110111011110001000011101100101001100100010001000100100011001100111011101110111011101110110011001100110010101010101010101000100010000110011001000100010001001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100101010101100111011101110110011001110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100101001100110011001101000100010001010101011001110111011101111000100010001000010100100010001000100011010101110110011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011000100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101000100010001000100010000110100001100110011001100110011001100110011001100110100010001000100010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110101011001100110011001100110010101100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100110011001000100011001100110011001100110101011101111000011110001000100001110110001100100010001000100101011101111000100001110111011101110111011101100110011001100110010101010101010001000100001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110010101100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100101001100110011001101000100010001010110011001110111011101111000100010001000011001000010001000100011010001110111011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010000100100010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001010100010001000100001100110100001100110011001100110011001100110011001100110100010001010101011001110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011101100110011001110110011001100110100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100010001100110011001101000111011101111000100010001000100010000110001000100010001001000110011110001000100010001000100010000111011101110111011101110110011001010101010001010100001100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110100001100110011001101000100010101010110011101110111011110001000100010001000011101010010001000100011010001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010000100100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001010101010101010101010001000100010000110011001100110011001100110011001101000100010101100111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001110110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001100110011010001100111011110001000100010001000100010000101001000100010001101010111100010001000100010001000100010001000011101110111011101110111011101100101010101010100001100100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100011001100110011001101000100010101010110011101110111100010001000100010001000100001100010001000100011010101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001010101010101010101010101100101010101010100010000110011001100110011010001000011010001000101010101100110011001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100011001100110011001000100010001000110011010001101000100010001000100010001000100010000101000100100010010101101000100010001000100010001000100010001000100001110111011101110111011101110110010101010100001100110010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100111100010000111011101111000011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000011001100110011010001000101010101100110011101111000100010001000100010001000100001100010001000100011010101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110010101000100010001000100010001000101010101010101010101000100001100110011001100110011010000110100010101010101011001100110011001100111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011101111000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000011001100110011001100110011001100110011010101101000100010001000100010001000100010000011001000100010011001111000100010001000100010001000100010001000100001111000100010001000011101110111011001010100001100110010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100111011110001000011110000111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010100110011001100110011010001000101010101100110011110001000100010001000100010001000100001110010001000100011010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100101010101010101010101010101010101100110011001100110011001010100001100110011001100110011001100110011010101010101011001100110011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010000110011001100110011001100110011001100110011010101101000100010001000100010001000100001110011001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010000111011001010100010000110010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010000111100001110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110010100110011001100110100010001000101011001100110011110001000100010001000100010001000100001110011001000100011010101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011001100110011001100110011001100110011001100110011001100101010001000100001100110011001100110011001100110011010001000101011001100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001100110011001100100011001100110011001100110011010001110111100010001000100010001000100001110011000100010011010101111000100010001000100010001000100010001000100010001000100010001000100010000111011001000101010000110011001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010000111100010000111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110010000110011001100110100010001000101011001100111011110001000100010001000100010001000100001110011001000100011010101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111010101000100010001000100001100110011001100110011001100110011001100110100010101100111011101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110011001111000011101100111011110001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100001010011001100110011001000100011001100110011001100110011010001110111011110001000100010001000100001100010000100010010011110001000100010001000100010001000100010001000100010001000100010001000100010000110010101100110010000110011001000100010001000110101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110010000110011001101000100010001010110011001110111011110001000100010001000100010001000100010000011001000100011010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110101010001000100010001000100001100110011001100110011001100110100001100110011010001000101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110011001111000011101100110010101100110010101010110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000100001100110011001100110011001100110011001101000100001101100111011110001000100010001000100101100010000100010011011110001000100010001000100010001000100010001000100010001000100010001000100001110101011001110101010001000011001100100010001000110011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110101010000110011010001000100010001010110011001110111100010001000100010001000100010001000100010000100001000100011011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101010100010001000100010001010100001100110011001100110011001100110100010001000011010001000100010001100111011110001000100010001000100010001000100010001000100010001000011110001000100010001000100001110111011001100110010101100111011001010101010101000100010001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010101010100001100110011001000100011001100110011001101000101010001010111011110001000100010001000100001010001000100100100100010001000100010001000100010001000100010001000100010001000100010001000011101100111011101100101010101010100001100100010001000110011010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110101001100110100010001000100010001010110011101110111100010001000100010001000100010001000100010000100001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110010000110100010001000100010101010100001100110011001100110011001100110011010001010100010001000100010001000101011110001000100010001000100010001000100010001000100010001000100001110111100010001000100001110110011001010110011001100110011001100101010001000100010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001000011001100110011001100110011001100110011010001000101010001000111100010001001100110001000100001000001001000100101100010001000100010001000100010001000100010001000100010001000100010001000011001111000011101100110010101010100010000100010001000110011010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110100001100110100010001000100010001010110011101110111100010001000100010001000100010001000100010000101001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100100010001000100010001000100010101010011001100110011001100110011001100110011010001010101010001000100010001000100010101100111100010001000100010001000100010001000100010001000100010000111011110001000100010000110010101010101011001010110011001010100010001000100010101010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010101000011001100110011001100110011001101000100010001000101010101010110100010001001100010001000100001000001000100100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100110010101010101010000100010001000110011010001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100100001101000100010001000100010101010110011101111000100010001000100010001000100010001000100010000101001000100011010101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101000100010001000100010001000100010101000011001100110011001100110011001100110011010001000101010101000100010001000100010101010110011110001000100010001000100010001000100010001000100010001000011001100111100010000111010101010101010101010101010101000100010001000100010001010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101010000110011001100110011001100110011001101000100010001000110010101010101011010001000100010001000100000110001000100100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001110110010101100101010000100010001000110011010001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010100010001000100010001000101010101100111011110001000100010001000100010001000100010001000100010000100001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110101010001000100010001010100010001000100010101000100001100110011001100110100001100110100010001000101011001010100010001000100010101010101011001111000100010001000100010001000100010001000100010001000100001100110011110000110010101010101010101010100010001000100010001000100010001010110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110100001100110011001100110011001100110011010001000100010001000110011101010110011001111000100010001000011100110001000100111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000110011001100101001100110010001000110011001101000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010100010001000100010001010101010101100111011110001000100010001000100010001000100010001000100010000100001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010100010001000100010101000100010001000100010001000100001100110011001101000100001100110100010001000101011001100101010001000101010101010101010101100111100010001000100010001000100010001000100010001000100001110110010101100111010101010101010001000100010001000100010001000100010101010110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010100001100110011001100110011001100110011010001000101010101000110100001110110011101111000100010001000011100100001000101001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000110011001100101001100110011001100110011001101000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010100010001000100010101010101010101100111011101111000100010001000100010001000100010001000100010000100001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101000100010001000100010001010101010001000100010001000100001100110011001101000100001101000100010001000100011001100110010101000101010101010101010101100111100010001000100010001000100010001000100010001000100010001000011001010101010101010100010001000100010001000100010001000100010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010011001100110011001100110011001100110011010001000101010101010101011110000110011110001000100010001000011000100001001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110101001100110011001100110011001101000101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001000100010001000101010101010101011001100111100001111000100010001000100010001000100010001000100010000101001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010000111011110001000011101110110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100001110101010001000100010001000100010101010101010001010100010001000100001100110011001101000100001101000100010001000100011001100110010101010101010101010101011001100111100010001000100010001000100010001000100010001000100010001000100001110101010001000100010001000100010001000100010001000101010101010110011101110111100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000011001100110011001100110011001100110011010001000110011001110110011110000111011110001000100010001000011000100001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110100001101000100001100110011001101000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101000101010001000101010101010101011001100111100010001000100010001000100010001000100010001000100010000101001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100111100010001000011001110111011101100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000011101010100010001000100010001010101010101010101010101010100010001000100001100110011001101010100001100110100010001000100010101100110011001100101010101010110011001100111011110001000100010001000100010001000100010001000100010001000100010000111011001010100010001000100010001000100010001000101010101010101010101100111011101111000011110001000011101100110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000010100110011001100110011001100110011001100110011010001010110011101110111011110001000011110001000100010001000010100100001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110100010001010100010000110011001101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010101010101010001010101010101100110011001100111100010001000100010001000100010001000100010001000100010000110001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000010010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110011110001000011101100110011101100110011001100111011101010110011110001000100010001000100010001000100010001000100010000111010001000100010001000100010101010101010101010101010101010100010001010100001100110011001101000100010001000100010001000100010101100111011101100110010101010110011001100111100010001000100010001000100010001000100010001000100010001000100010001000011001010100010001000100010001000100010001000101010001000101010101100111011101110111011101110111011001100110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010000110011001100110011001100110011001100110011010001010110011101110111100010001000100010001000100010001000010100100001001001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100100011001100101010101000011001101010110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010101010101010001010101010101100110011101110111100010001000100010001000100010001000100010001000100010000110001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000110101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100101010101100111011101110101010101100110010101010111011101010110011110001000100010001000100010001000100010001000100001110101010101010100010001010101011001100110011001100110011001010101010101010100001100110011001100110011010001000100010001000100010101100111011101100110011001100110011001111000100010001000100010001000100010001000100010001000100010001000100010000110010101000100010001000011001100110011001101000100010001000101011001110111011001100110011001100110011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100101110100010000110011001100110011001100110011001100110100010101010110100001111000100010001000100010001000100010001000010100100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100101011101100101010100110011010001010111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101010101010101010101010101100110011101110111100010001000100010001000100010001000100010001000100010000111001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001100110011001010101011001100110010101010101010101010110011001010110011101110111011110001000100010001000011101110111011101110111011001010101010101010101011001100110011001100110011001010101011001010100001100110011001100110011001100110100010001000101010101010111011101110110011001100110011001111000100010001000100010001000100010001000100010001000011110000111100001110101010001000100010001000011001100110011001100110100010001000101011001100110011001100110011001100110011001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010100010100110011001100110100010001000100001100110100010101100110100010001000100010001000100010001000100010001000010000100001001110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010110011101100110010100110011010001010111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010101010101010101100101010101100110011110001000100010001000100010001000100010001000100010001000100010000111001100100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110110011001100101010101010101010101010101010101010100010101010101010101010110011001100111011110001000100010000111011001100110011101110111010101010101011001010101011001100110011001110111011001100110011001010100001100110011001101000100010001000100010001000101010101010110011101110111011101110110011001111000100010001000100010001000100001110111011001100110010101010101010101010110010101000100010001000011001100110011001100110100010001010101011001100110010101100110011001100110011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001010110011001000011010001000100010001010101010001000101011001100111100010001000100010001000100010001000100010000111010000100001010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100111011101100110010000110011001101010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101010110010101100101011001110111011110001000100010001000100010001000100010001000100010001000100010001000001100100010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001110110011001010101010101010110010101010101010101010100010001000100010001010101011001100111100010001000011101100110011001110111011101110110010101100110011001010110011001100110011001110111011001100110011001010100001100110011010001000100010001000100010001000101010101010110011101110111011101110110011001111000100010001000100010001000011101110110011001100110010101010100010001000100010001000100010000110011001100110011001100110100010101010101010101010101010101100110011001100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100111010100110100010001000100010001010110010101010110011001110111100010001000100010001000100010001000100010000111001100100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001110111011101100110010000110010001101010111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101100110010101100110011001110111011110001000100010001000100010001000100010001000100010001000100010001000010000100010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100001010010000100100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011001100110010101010101010101010110011001010101010101000100010001000100010001010101011001100111100010001000011001100101011001110111011101110111011101110110011001100111011101110110011101110111011001100110010101000100010001000100010001000100010001000100010001010101011001010110011101110111011101110111011001111000100010001000100010000111011101100111011101110111011001010101010001000011001101000100010001000011001100110011001101000100010101010100010001000100010101010110011001100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001110110010001000100010101010101010101100111011001100110011101110111100010001000100010001000100010001000100010000111001100100001010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110010000110010001101010110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100110011001100110011101110111011110001000100010001000100010001000100010001000100010001000100010001000010000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000100001000001000100100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110010101010101010101000101011001100101010101000100010001000100010001000101011001100111011101110110011001010110011101110111011110000111011101100110011001110111011101110110011101110110011001110110010101000100010001000100010001010100010001000100010101010110011001100110011110001000011101110111011001111000100010001000100010000111011101111000100010000111011001010101010001000100001100110011010001000011001100110011001101000101010101000100010001000100010101100110011001100111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001010101010101000100010101010110010101100111011110000111011110001000100010001000100010001000100010001000100010000110001100100001010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111011001100101010100110010001101000110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100111011001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000010100100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000011100110001001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011001010101010001000100010001010110010101000100010001000100010001000101011001110111011101100110010101100111011101111000100010000111011101110111011101110111011101100110011101110110011101110110010101010100010001000100010101010101010001000101010101010110011001110110011110001000100001110111011101111000100010001000100010001000100010001000100010000111011001010100010001000100001100110011001100110011001100110011001100110100010001000100010001000100010101010101011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101010101010101000100010101100111011001100111100010000111011110001000100010001000100010001000100010001000100010000110001100100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101100110010100110010001001000110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000011000100001000100100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001010101010001000100010001000100010101010100010001000100010001000101011001100111011001100101011001100110011101111000100010001000011101110111011101110111011101100110011101100110011101110110010101010100010001000100010101010101010101010101010101010110011101110110011110001000100010001000011101111000100010001000100010001000100010001000100010000110011001010100010001000100001100110011001100110011001100110011001100110100001100110100010001000100010001000101011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010101010101010101000101010101100111011101110111100010001000011101111000100010001000100010001000100010001000100010000110001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001110111011000110010001000110110011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001100111011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000011000100001001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110110010101010101010001000100010001000100010001010100010001000100010001000101011001100101010101010101010101100110011101111000100010001000100010000111011101110111011101100111011101100110011101110110010101010100010001000100010101010101010101010101010101010110011101110111011010001000100010001000100001111000100010001000100010001000100010001000100001110110011001010101010001000100001100110011001100110011001100110011001100110100001100110100010001000100010001000101011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110101010101010101010101010101011001100111011101110111100010001000011110001000100010001000100010001000100010001000100010000110001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010110100010000111011000110011001000110101011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010001000001100010001001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101100110011001100110010101010100010001000100010001000100010001000100010001000101010101010101010101010101011001100110011101111000100010001000100010001000100001110111011001100110011101010110011001100110010101000100010001000101010101010101010101010101010101010101011001110111011010001000100010001000100010001000100010001000100010001000100010001000100001110110011001010101010001000100001100110011001100110011001100110011001101000100001100110100010001000100010001000100010101010101011001100111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100101010101010110010101010101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101101000100010001000011000110011001000110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010000111001100010001001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110110011001100110011001100110011001100101010101000100010001000100010000110011001101000100010001000100010101010100010001010110011001100111011101111000100010001000100010001000100001110111011001010101010101010101010101010101010101000100010001000101010101010101010101010101010101010101010101110111011010001000100010001000100010001000100010001000100010001000100010001000011101110110011001010100010001000100001100110011001101000100001100110011001101000100010000110100010001000100010001000100010101010110011101110111011101111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110010101010110010101010110011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000011000110011001100110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010000110001000010001001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101100101010101010101010101010100010001000100010001000100001100110011001101000100010001000100010001000100010101010111011101110110011001110111100010001000100010001000100001100101010101010100010101010101010101010101010101000100010001010101010101100101010101010101010101010101011001100111011001111000100010001000100010001000100010001000100010001000100010001000100001110110011001100101010001000100010001000100010001000100010000110011001100110100010001000100010001000100010001010110011001110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100110010101100110011001100110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000110011001100110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100000110010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100010000100001000010001001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100101010101010101010101010100010001000100010000110011001100110100001101000100010001000100010001000100010101100111011001110111011101110111100010001000100010000111011001010101010101010101010101010101010101010101010101000100010001010101010101100110011001010101010101010101011001100110011001111000100010001000100010001000100010001000100010001000100010001000100001110111011101100101010001000100010001000101010101010101010100110011001100110100010001000100010001010101010101100111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110011001100110011001110110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000110011001100110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100000110001001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100001110011001000010001001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001100110011001100101010101000100010001000011001100110011001100110100001101000100010001000100010001000101010101100110011001100110011101110111100010001000100001110110010101010101010101010101010101010101011001100101010101000100010001010101010101100110011001100101010101010101011001100110011001111000100010001000100010001000100010001000100010001000100010001000100001110111011101100110010101000100010001000101010101100101010000110011001100110100010001000100010101010101011001100110011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110011001110110011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000011001100110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000001001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100001110010000100010010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100110011001010101010101000100010001000100001100110011001100110011001100110100010001000100010001000101011001100110011001100111011101111000100010000111011101100110011001100101010101010101010101010101010101010101010101000100010001010101010101100110011001100110011001010101011001100111011001111000100010001000100010001000100010001000100010001000100010001000100001111000011101110110010001000100010001000101011001100100001100110011010001000100010001000100010101100110011001100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101100111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000011001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000100001100110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100001010010000100010010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100101010101000100010001000100001100110011001100110011001100110011001100110100010001010101011001100110011001100111011101111000100001110111011101100110011001010101010101010101010101010101010101010101010101000100010101010101011001100110011101100110011001100101011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000011101100100010001000100010001010110011001000011001100110011010101100101011001010100010101010110011001100110011001100111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001000100001101000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000100001000010000100010010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011001100101010101000100010001000100001100110011001100110100001100110011001100110100010001010110011001100101011001100111100001110111011101110111011101100101010101010101010101010101010101010101010101010101010101000100010101100101011001100110011101110110011001100110011001100111011110001000100010001000100010001000100010001000100010001000100010001000100001110110010101000100010001000101010101100110010000110011001100110011001101010110011001100110010101010101010101010110011101110111011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000100001101000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000011100110001000100100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100101010001000100010001000011001100110011001100110011001100110011001100110100010101100110011001010101011001110110011001010101010101010110011001100101010101010101010101010110010101010101010101010101010101000100010101100110011001100111011101110111011101100110011001100111011110001000100010001000100010001000100010001000100010001000100010000111010101010100010001000100010001010110011001100101001100110011001100110011001101000100010001000100010001010110010101010101010101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010101010001000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000011000100001000100100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001010101010101010100010000110011001100110011001100110011001100110011010001000100010101010101010101010101010101000100010001010101010001000101011001100101010101010101010101010101011001010101010101100101010101000101010101100110011001110111011101110111011101110111011001111000100010001000100010001000100010001000100010001000100010001000011101100101010001000100010001000101010101100111011001010011001100110011001100110011001100110011001101000100010001000100010101100101010101010110011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010101010001000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010001000010000100001000100100010010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110010101010101010101000100010000110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010101100110011001010101010101010101010101100101010101010101011001100101010101100101010101000101010101100110011001110111011101110111011101110111011001110111100010001000100010001000100010001000100010001000100010000110010101000101010101000100010001010101011001100110011001000011001100110011001100110011001100110011001101000100010001000100010001010110011001010101010101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100011001000010100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100110010001000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110010001000100010001110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010000111001100010001000100100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100101011001100110010101000100010000110011001100110011001100110011001100110011001100110011010000110011001101000100010001000100010101110111011101100110010101010101010101100110011001010110011001100110010101100101010101010101010101100110011001110111011110001000100001110111011001110111100010001000100010001000100010001000100010001000011001010101010101010101010101010101010101010110011101100110010100110011001100110011001100110011001100110011001101000100010001000100010101010101010101100110010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101100110010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110010000100100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010000110001000010001000100100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001100110011101110110010101000100010000110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010101100111011101110111011001010101010101010110011001010110011001100110010101010101010101000101011001100110011001110111100010001000100001110111011110001000100010001000100010001000100010001000100001100101010101010101010101010101010101010101011001100111011101100110010000110011010000110011001100110011001100110011001100110100010001000100010001010101010101100110011001010101010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110010101010110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011000100010010001001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100010000101000100010001000100100101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001111000011101100101010101000100010000110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010101100111011101110111011101100101010101010101011001010101011001010110011001010101010101010101010101100110011101111000100010001000100010000111011110001000100010001000100010001000100010000111011001010101010101010101010101010101010101010110011101110111011101100101010000110011001100110011001100110011001100110100010001000100010001000101010001010101010101100110011001100101010101000101011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011000100010010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100001110011000100010001001000110110011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110110010101000100010001000011001100110011001100110011001100110011001100110011001100110011010001000100010001010101010101100111011101110111011101110110011001010101010101010101010101010110011001100100010101010101010101100110011101111000100010001000100010001000100010001000100010001000100010001000100001100110010101010101010101010101010101010101010101100111011101110111011101100100010001000011001100110011001100110011001100110100010001000100010001000101010101010101011001010101010101010110010101010101011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000011000100010010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100001100010000100010001001000110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100001110111011001010100010001000011001100110011001100110011001100110011001100110011001101000100010001000101010101010110011001100111011101110111011101110111011001100101010101010101010101010111011101100100010001010101010101100111011101111000100010001000100010001000100010001000100010001000100010000111011001010101010101010101010101010101010101010101011001110111011101110111011001000100010001000011001100110011001100110011001100110100010001000100010001010101010101010101010101010101010101010110011001100101010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100000100100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000100001010010000100010001001001000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011101110111011101010100010001000100010001000100001100110011001100110011001100110011010001000101010101000100010001010101010101010110011101110111011101110111011001100101010101010101010101100110011001010100010001010101011001100111011110001000100010001000100010001000100010001000100010001000100001110101010101010101010101010101010101010101010101010110011001110111011101110111010100110100010001000011001100110011001100110011001100110011010001000100010101010101010101010101010101010101010101010110011001100110011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000011101000001000100010001001001010111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011001100110010101010101010101010101010101010101011001110111011101100100010001000100010001000100010000110011001100110011001100110011001101000100010001000100010001000100010001000101011001110111011101110111011001100110011001010101011001100110011001010100010001010101011001100111100010001000100010001000100010001000100010001000100010001000011101010101010101010101010101010101010101100101011001100111011101110111011101110111010001000100010000110011001100110011001100110011001100110011001101000100010101010101010101010101010101010101010101010110011001100110011001100110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000011000100001000100010010001101101000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000011101110110011001010101010101010101010001000101010001000100010001000100010000110011010001000100010101010100010001000101010101010101010001000011001100110011001100110011001100110011001100110011010001000011010001000100010001000101011001100111011101110110011001010101011001100110011001010100010101010101011001110111100010001000100010001000100010001000100010001000100010000111010101010101010101010101010101010101010101010110011001110111011101110111011101110101010001000100010000110011001100110011001100110011001100110011010001000100010001010101010101010101010101010101010101010110011001010110011101110111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010001000010100100001000100010010010001111000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010000111011001010101010101010101010101010100010001000101010001000100010001000100010001000100010001000100010000110011001100110011001100110011010001000100010001000011001100110011001100110011001100110011001100110011001100110011010001000100001101000100010101010110011101110111011101100101011001100110011001010100010001000101011001110111100010001000100010001000100010001000100010001000100001110110010101010101010101010101010101010110010101100111011101110111011101110111011101000100010001000100010000110011001100110011001100110011001101000100010001000100010001000101010101010101010101010101010101010110011001010110011101110111011101110110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010000111010000010001000100010010010001111000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010000111011001010101010101010101010101010101010001000100010001010101010101010101010001000101010101010100010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010000110011001101000100010001000100010101010101010101100111011101100101011001100110011001000100010001010101011001111000100010001000100010001000100010001000100010001000011101100101010101010101010101010101011001100101010101110111011101110111100010000110010101000100010101010100010000110011001100110011001100110011001101000100001100110100010001000101010101010110010101010101010101010110011001100110011001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010000111001100010001000100010010010110001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000011101100101010101010101010101100110010101010101010101010101010101010110011001100110010101100110011001100101010001000100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000101010101010101010101010111011101100110011001100110011001000100010101010110011101111000100010001000100010001000100010001000100010001000011101100101010101010101010101010110011001100101011001110111011101110111011101100101010001010101010101010100010001000100001100110011001100110011010001010100010000110100010001000100010101010101010101010101010101010110011001100110011001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010000110001000010001000100010011011010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010000111011001100110011001100110011001100110011001010110011001100110011001100111011101100110010101100111011101100101010101010101010101010100001100110011001100110011010001000100001100110011001100110011001100110011001100110011001100110100010001000100010101010101010101010110011001100110010101010110011101110110011101110111011001000100010101010110011110001000100010001000100010001000100010001000100010001000011001100101010101010101011001100110011001110110011101110111011101110101010001000101010101010101010101000100010001000011001100110011001100110011010001010100010001000100010001000100010001010101010101010101010101010101011001100110010101100111011110000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100010000100001000010001000100100011011110001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100001110110011001100110011001100110011001100110011001100111011101110111011101110111011101110110010101110111011101110110011001100110010101000011001100110011001101000100010001000011001100110011001100110011001100110011001100110011001101000100010001000011001101000100010001000101011001100110011001100110011101100101011001100111010101000100010101010111100010001000100010001000100010001000100010001000100010000111011001010110010101100110011001100111011101110110011110000111010101000101010101010101010101010101010101000100001101000011001100110011001100110011010101010100010001000100010001000100010001010101010101100110010101010101011001100110011001100111100010000111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100001110011000100010001000100100100011110001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100001111000011101100111011001100110011001110111011101110111011101110111011101110111011101110111011101110110011101110111011101110110011001100101010000110011001100110100010001000100010001000011001100110011001100110011001100110011001100110011010001000100010000110011001100110011001100110100010001010110011001100110011101010100010101100111010101000100010101100111100010001000100010001000100010001000100010001000100010000111011001100110011001100110011001110111011101110111011101110101010101010101010101010101010101100110010101000100010000110011001100110011001100110011011001010100010001000100010001000100010001000101011001100110010101100110011001110111011001100111100010001000011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100001100010000100010001000100100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100111100010001000011101111000011101100111011001100111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100110011001010011001100110011001100110100010001010101010000110011001100110011001100110011001100110011001100110011001101000101010001000011001100110011001100110011001101000100010001010110010101000100011001110110010001000101010101100111100010001000100010001000100010001000100010001000100010000111011001100110011001100110011101110111011101110111011001010101010101010101010101010101011001100110010101000101010001000011001101000011001100110011010001000100010001000011001101000100010001000100010101100110011001100110011001100111011001100111100010001000100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100001100010000100010010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101101000100010001000100010000111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101100110010000110011001100110011001101000100010001010101001100110011001100110011001100110011001100110011001100110011001100110100010101010100010000110011001100110011001100110011001101000100010001000100010101110110010001000100010101101000100010001000100010001000100010001000100010001000100010000111011001110111011101110111011101110111011101110111010101010101010101010101010101010101011001110110010001000101010001000011010000110011001100110011010001000100010001000100001101000100010001000100010001010110011001100110011001100110011001100110100010001000011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000100011100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000100001000010000100010010001001000111100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100001110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010100001100110011001101000100010001000100010101010100001100110011001100110011001100110011001100110011001100110011001100110100010001000101010000110011001100110011001100110011001100110011001101000100010101100101010001010101010101111000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110101010001010101010101010101010101100110011101110101010001010101010000110100010000110100001100110011010001000100010001000100010001000100010001000100010001000101011001100110011001100111011001100110011110001000011101100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000011100110001000100010010001001011000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001000100010000110011001101000101010001000101010101000011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000011001100110011001100110011001100110011001100110100010001100101010001000101011001111000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010100010001010101011001100111011101110100010001100101010001000100010000110011001100110100010001000100010001000100010001000100010001010100010001000100010101100110011001110111011101100110011110001000011001100110011110001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100000110010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000011000100001000100010010001001101000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010000110011001100110011010001010100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000011001100110011001100110011001100110011001100110100010001010100010001000101011001111000100010001000011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101000100010101010110011001110111011101010100010101010100010001000100010000110011001100110100010001000100010001000100010001000100010001010101010101010101010101010110011001100111011101100110011010000111010101010110011101100101010101100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010001000010000100001000100010010001101111000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100001100110011001100110011001101000100010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100001100110011001100110011001100110011001100110011010001000100010001000101011010001000100001110110010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010001000100010101100110011110001000011101000100010001000100010001000100010000110011010001000100010001000100010001000100010001000100010001010110010101010101010101010110011001100111011101100110011010000110010001010101010101010101011001100111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010000111001100010001000100010010010010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010001000100001100110100001100110011001101000101010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010000110011001100110011001100110011001100110011010001000100010001010101011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000100010101000100010101100110011110001000011001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001010101010101010101010101010101011001100110011101100110011001110110010001010100010001010101011001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010000110001000010001000100010010010110001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000100010001000100001100110100001100110011001101000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011001100110011001100110011001100110011001100110100010001000101011001100110010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010001000101010101000100010101100111011110000111010101000100010001000100010001000100001100110100010001000100010001000100010001000100010101000100010001010101010101010101010101010101010101100111011101110101010101100101010101010100010001010101011001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010000101001000010001000100010010011010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001000100010001000100010001000100010001000100010001000011110000110011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100010001000100001100110100001100110011010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010100010001010101010101100111011110000110010001000100010001000100010001000100001100110011010001000100010001000100010001000100010101010100010001010101010101010101010101010100010101100111011101110101010001010100010101010100010001010110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010000100110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100010000011000100010001000100100011011110001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100100010001000101010101000100001101000100001100110100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101100100010101000100010001010110011001100111011101110101010001000100010001000100010001000100010001000100010001000100010001000101010001000101010101010100010001010101010101010101011001100101010101010110011101100101010001010100010001000100010101100110011101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100001100010000100010010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100001110110011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101111000011101010101010101010101010101000100010001000011001100110100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000011010001000100010001010101011001110111011101110111011101110111011101110111011001110111011101110111011101010100010001000100010001010110011101110111011101110100010001000100010001000100010001000100010001000100010001000100010001010101010101010101011001100100010101100110010101010101011001100110010101010110011001110110010001000100010001000101011001100111011101110111011101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100001010010000100010001000100100110100010001000100010001000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011110000111011001010101011001100110010101000100010001000100001101000100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001010101010101100110011001100110010101100110011001100110011001110111011101110111011101010100010001000100010001010101011001110111100001110100010001010100010001000100010001000100010001000100010001000100010101100101010101010110011001100101010001100111011001100101010101010101010101010101011001110110010001000100010001000101011001110111011101110111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000100000110001000100010001000100110111100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010001000100010001000100010001000100010001000100001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110000110010101010101011001100110010001000100010001000100001101000100010101000100010000110011001100110011001100110011001100110011010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010101010110011001100110010101100110011101110111011101110111011101110111011101000101010101000100010001010110011101110111011101100100010101010101010101000100010001000100010001000100010101000100010101100101010101010110011001100101010101110111011001110110011001010101010101100110011001100101010001000100010001010110011001110110011001100110011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000011100100001000100010001000101001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011010001000100010001000100010001000100010001000100010001000100010001000100001100111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011101110111100001110101010101010101011001100110010001000100010001000100010001000100010101000101010000110011001100110011001100110011010000110011010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000101010101010101010101010101011001100110011001100110011001110111011101110111011001000101010101000101010101010110011101110111011101010100010101010101010101010101010101000100010001000100010001000100010101100101011001100111011101110110010101110111011101110111011001100101010101010110011001010100010001000100010001100110011001100110010101010101011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000010100100001000100010001000101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011010001000100010001000100010001000100010001000100010001000100010001000011101100111011101110111011101110111011101110111011101110111011101110111011101111000011101111000011101110111011101100101011001100110011001100101010001000100010001000100010001000101010101010101010000110011001100110011001100110011001101000100010000110011001100110100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001010101010101010101010101100110011001100111011101110111011101110111011101110111010101000101010101000101010101010111011101110111011101000101011001010101010101010101010001000100010001000100010001000100010101010110011001100111011101110110010101100111011101110111011001100110011001010101010101010100010001000100010101100101010101010101010101100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000010010001001000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010001000001100010001000100010001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000100010001000100010001000100010001000100010001000100010001000011101010111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101111000011101010101010101010110011001100101010001000100010001000100010001000101011001100101010000110011001100110011001100110011010001000100010001000011001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001010101011001010100010101010101011001100110011001110111011101110111011101110111010101000101010101000110011001100111011101110111011000110101011001100101010101010101010001000100010001000100010001000101010101010110011001100110011101110110010101100111011101110111011101100110011001100101010101000100010001000100010101010101010101010101010101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010000111001000010001000100010001001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001111000100010000111100010001000100010001000100010001000100001111000011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010101010110011001100101010001000100010001000100010001000101011101100100010000110100001100110011001100110011010001000101010001000011001101010100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000101010101010100010001010100010001010101011001100110011001100111011101110111011101110111011001000110011001010110011001100111011101110111011001000110011001100101011001010101010001000100010001000100010001000101011001010111011101110111011101100110010101010110011001100110011001110110011001100110010101010100010001000100010101010101010101010101010101010101011001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010000100110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010000101001000010001000100010001010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001101000100010001000100010001000100010001000100010001000100010001000011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101010101010101100110011101100101010001000100010001000100010001010101011101100100010001000100001100110011001100110011010101010101010100110011001101010100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011010001000100010001000100010001010101010101100110011001100111011101110111011101110111011001000110011001010111011101110111011101111000010101000111011001100110011001100110010101000100010001000100010001000101011001010110011101110111011101100110010101010101010101010101010101100101010101010100010001000100010001000100010001010101011001100110011001100110011001100110011001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100010000100000100010001000100010001010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101101000100010001000100001111000100010001000100010001000100010001000010101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110110010101010101010101010110011101100100010001000100010001000100010001010110011001010100010001000100010000110011001100110011010001100110010000110011010001010101010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001010101011001100110011001100111011101110111011101110111011001000110011001100111011101110111011101110111010001010111011001100111011001100110010001000100010001000100010001000110011001000110011101110110011001110110010101010101010101010101010101010101010101010100010001000100010001000100010001010110011001100110011001100111011101110111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100001110010000100010001000100010010011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101101000100010001000100010001000100010001000100010001000100010000111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010101010101010101011001010100010001000100010001000100010001010110011101010101010001000100010000110011001100110011001100110100001100110011010001010110010001000011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000101010101100110011001110111011101110111011101110111011001010110011001100111011101110111011101110111010001100111011101110111011101110110010101010100010001000100010001010110010101000110011101110110010101010101010101010101010101010101010101100101010001000100010001000100010001000100010001000101011001100110011001100111011101110111011101110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100001010010000100010001000100010100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101010111100010001000100010001000100010001000100010001000100010000111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101010101010101010101011001010110010001000100010001000100010001010101010101010111011101010100010001000100010000110011001100110011001100110011001100110011001101000101010000110011001100110011001100110011001100110011001100110011001000100011001100110011001100110011001100110011001100110011001100110011001100110011010001000100001101000100010001000101010101100110011101110111011101110111011001010110011101100111011101110111011101110110010001100111011101110111011101110111011001010100010001000100010001010110010101000110011001100111011101100101010101010110011001100110011001010100010001000100010001000100010001000100010001000100010001000101011001100110011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000100001000001000100010001000100010101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100111100010001000100010001000100010001000100010001000100010000110010110000111100001110111011101110111011101110111011101110111011101110111100010000111011101110111010101010101011001100110010101010101010001000100010001000100010001010101010101100111011101100101010001000100010001000100010000110011001100110011010101000011001101000101010101000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010000110011001100110011001100110011001100110011001101000100010001000100010001000100010101010110011001110111011001010110011101100111011101110111011101110110010001110111011101110111011101110111010101010100010001000100010001100110010101010110010101100110011001010101010101010110011001100111011001000100010001000100010001000100010001000100010001000100010001000100010101010101011001100111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000011000100001000100010001000100100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100111100010001000100010001000100010001000100010001000100010000110011010000111100010000111011101110111011101110111100001110111011101110111011101110111011110000111011001010101011101110110010101010100010001000100010001000100010101100101011001110111011101100101010001000100010001000100010000110011010001000100010101000011010001000101010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010000110100010001000100010001000101011001100111011001010110011101100111011101110111011101110101010101110111011101110111011101110110011001010100010001000100010001100111010101010110011001100110011001100110010101010101011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000100010011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000010100100001000100010001000101001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000100010001000100010001000100010001000100010000101011010000111011101110111011101110111011101110111011101110111011101110111011101111000100010000110010101010111011101110101010101010100010001000100010001000100010101100110011001110111011101100101010001000100010001010101010001000011010001010100010100110100010001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000101011001110110011001010110011101110111011101110111011101110100010101110111011101110111011101100110011001010100010001000100010001100110010001010110011001100101011001100110010101010110011101010100010001000100010000110100010001000100010001000100010001000100010001000100010001000100010101010101011001110111011101111000011101110111011101110111100001111000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010001000001100010001000100010001000101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110100010001000100010001000100010001000100010001000100001110101011101110111011101110111100001110111011101110111011101110111011101111000011101111000100010000111011001110111011101010101010101010100010001000100010101010101010101100111011001110111011101100101010101010101010101010101010100110011010101000100001100110100001100110011010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010101000101011001100111011001100110011101110111011101110111011101110100011001110111011101110111011101110111011001010100010101000100010101110110010001010110011001100110011001110110010101100110010101000100010001000100001100110011010001000100010001000100010001000100010001000100010001010101010101010101010101010111011101110111100001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010000110001000010001000100010001001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110100010001000100010001000100010001000100010001000100001110101011110000111100001111000100001110111011101110111011110000111011101110111011110001000100010000111011101110111011001010101010101010100010001000100010101010110011001100111011101110111011101110101011001010110010101100101010000110011010000110011001100110011001100110100010101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010101010101010101010101010101100110011001100110011101110111011101110111011101100100011101110111011101110111011101110111011001010101010101000100010101110110010001010110011001100110011101110110011001100101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101011001010101011001010101011001110111011101111000100001110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100010000101000100010001000100010001001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110110100010001000100010001000100010001000100010001000100001110101100010001000100001110111011101110111011101110111011110001000100010000111100010001000100010000111011101100110011001100101010101000100010001000101010101100111011101110111011101110111011101110110011001100110011001100101001100110011001100110011001100110011001101000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010000110100010001000101010101010101011001100110011001110110010101110111011001100110011101110111011101110111011101010100011101110111011101110111011101110111011001010101010001000100011010000110010001100110011001100110011101110110011101010100010001000011001101000100010001000100010001000100010001000100010001000100010001000100010001000101011001100110010101100101010101100111011101111000011101110111011110001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100001110011000100010001000100010001010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011110001000100010001000100010001000100010001000100001100101100010001000100001111000100001110111011101110111011110001000011101111000100001111000100001110110011001101000011101010101010101000100010001000101011001110111011101110111011101110111011101110110011001100111011001010011001100110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001010101010101010101010101010100010001000100011001100110011101110111011101110111011101100110011101110111011101110111011101110111011101010101011101110111011101110111011101110111011001010101010001000100011110000110010001100110011001110111011101110111010101000100010001000011010001000100010001000100010001000100010001000100010001000100010001010100010001000101011001100110011001100110011001010110011101110111011101110111011101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100001100001000100010001000100010001011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101011110001000100010001000100010001000100010001000100001010110100010001000100010001000100010000111011101111000100001110111011101111000100010001000100001110101011010001000011001010101010101010100010001000101011001110111011101110111011101110111011101110111011101110111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001100110010001100110011001100110011001100110011010001000100010101010110011001010101011001100101010001000110011101110111011101110111011101110110011001100111011101110111011101110111011101000110011101110111011101110111011101110111011001100110010001000101011110000101010001100111011101110111011101110101010001000100010001000100010001000100010001010100010001000100010001000100010001010101010001010100010001000100010101100111011101110110011001100110011001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100001000001000100010001001000010011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011010001000100010001000100010001000100010001000100001010111100010001000100010001000100001110111011101110111100001111000100010001000100010001000100001110111011110000111011001010101010101010101010001000101011101110111011101110111011101110111011101110111011101110101010000110011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110010001000110011001100100011001100110010001100110011001100110011010000110011001100110100010001000101010101010100010101010101010101000100010101010110011101110111011101110111011101100111011101110111011101110111011001000111011101110111011101110111011101110111011001100110010001000110011110000101010001100111011101110111011101100101010001000100010001000100010001000100010101010100010001000100010001000100010001010101010001000101010101010100010001010111011101110111011001100110011001101000011101110111011101110111011101110111011110001000011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001101010101010101010101001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b100000100001000100010001001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110011010001000100010001000100010001000100010001000011101000111100010001000100010001000100001111000100001111000011101111000100010001000100010001000100010001000100010000110011001010110011001100101010101010101011101110111011101110111011101110111011101110111011101100100001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100011001100110011001100110011001100110011001100110011010000110011001100110011001101000100010001000100010001010100010001010100010001000101011001100111011101110111011101110111011101110111011101110111010101010111011101110111011101110111011101110111011101110101010001000111011101110101010101110111011101110111011101100101010001000100010001000100010001000101010101000100010001000100010001000100010001010110010101000101010101010101010001000110011101110111011101100110011001100111011101110111011101110111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101010101010101010101010100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b010100100001000100010001000101001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110010110001000100010001000100010001000100010001000011001000111100010001000100010001000100001110111011101111000011110001000100010001000100010001000100010000111100001110101010101100111011001100110010101100101011101110111011101110111011101110111011101110111011001000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000110011001100110010001000110011001100110011001100110011001100110100010001000100001101000100010001000100010101000100010001000100010001000101010101010110011101110111011101110111011101110111011101110111010001100111011101110111011101110111011101110111011101110101010001010111011101110100010101110111011101110111011001100101010001000100010001010100010001010101010001000100010001000100010001000100010001000110011001000101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001101010101010101010101010101010101010101010101010101010011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100010001000100010001000101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010110001000100010001000100010001000100010001000011001011000100010001000011101111000100001110111011110001000011110001000100010001000011101111000100010001000100001100101010101110111011001100110011001110110011001110111011101110111011101110111011101110111011001010100001100110011001100110011001100110011001100110011001100100010001100100011001100110011001100110011001100110010001000100011001100110010001100110011001100110011001100110011001100110100010001000100001101000100010001000100010101010101010101000100010001000101010101010110011001110111011101110111011101110111011101110110010001110111011101110111011101110111011101110111011101110100010001100111011101110100010101110111011101110111011101100101010001000100010101010101010101010100010001000100010001000101010101000100010001000101011001010101011001100101010101010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011010101010101010101010101010101010101010101010101010101010011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001000110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001000100010001001001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010001111000100010001000100010001000100010001000010101101000100010000111011101110111011101110111011101110111100010000111011101111000011110001000100010000111011101100110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001100110010001000110011001100110011001100110011001100110011010001000100001101000100010001000101010001000101010101010100010001000100010001010101010101100111011101110111011101110111011101110101010001110111011101110111011101110111011101110111011101110100010001100111011101100100011001110111011101110111011101100101010101000101010101010101010101000100010001000100010001000101010101010101010001000100010101010101011001100110011001100101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001000100010010001110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010001101000100010001000100010001000100010000111010101101000100010000111100001110111011101110111011110001000100010000111011101110111011101111000100010000111011001100111011101110111011101100111011101110111011101110111011101110111011101110111011101110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000100010001100100010001100110011001100110011001100110011001100110011001100110100010001000100010001000101010101000101010101100101010001000101010101010101010101010110011001110111011101110111011101110100010101110111011101110111011101110111011101110111011101100100010101110111011101100100011101110111011101110111011101100110010101010110010101010101010001000100010001010100010001010101010101010101010001000100010101100110011001110111011101100110011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100011001000100011001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001000100100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101101000100010001000100010001000100010000111010001111000011110000111100001110111011110001000011110001000100010001000100010000111011110001000011110000111011001111000011101110111011101110111011101110111011101110111011101110111011101110111011101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000100011001100100010001000100010001100110011001100110011001100110011001100110011001100110100010001000100010001000100010101010101010101100110010101000101010101010101011001010101010101100111011101110111011101110011011001110111011101110111011101110111011101110111011101010100011001110111011101010101011101110111011101110111011101110110010101100110010101010101010001000100010001010101010001100110010101010101010101000100010001100110010101111000011101110110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101010101011101110111010101010111011101010101010101010101001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100011001100100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001000100100010011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010101011000100010001000100010001000100010000110010101111000100010000111100001110111011110000111011110001000100010001000100010000111011101110111011110000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111010100110100001100110011001100100010001100110011001100110011001100110011001100110011001100110011001100100010001000100010001000100010001100110010001000110010001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000101011001010101011001010101011001100110011001100110010101100110011001110111011101010011011101110111011101110111011101110111011101110111011101000100011101110111011101010101011101110111011101110111011101110111011001110111011001100101010001000100010001010101010101100110011001010101010101000100010001010110011001100111011101110110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101010111011101110111011101110111011101010101010101010101010100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100011001100100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001001000100100100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010000111011001100111010101101000100010001000100010001000100010000110010110000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001000100001100110011001100110011001100110011001100110011001100110011001101000100001100110011001100100010001000100010001000100010001100110010001000100010001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010101100101011001100101011001100110011101110110011001100110011001100111100001000100011101110111011101110111011101110111011101110111011101000101011101110111011101000101011101110111011101110111011101110111011001110111011101100101010001000100010101010101010101100110010101100110010101010100010001010111011001100111011101110111011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101110111011101110111100110010111010101111001100101110101010100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010010001000100110011101111000100010001000100010001000100010001000100010001000100010001000010101000101011001111000100010001000011101000011001100110101011001101000100010001000100010001000100010000101011010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001000100010001000100010001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000101011001110110011001110111011101110111011001110110011001100110011000110110011101110111011101110111011101110111011101110111011001000110011101110111011101000110011101110111011101110111011101110111011001100111011101010101010101010101010101010101010101100110011001100110010101010101010001010110011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101110111100110010111011110010111011110011011101110110111010100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001100100011001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001000100110101010001001000100010000111011010001000100010001000100010001000100010000110010001000100001101000101011001111000011100110011010000110100010001011000100010001000100010001000100001110100011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000100010001000100010001000100010001100110010001000110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010101100110011001110111011101110111011101110111011001100110010100110111011101110111011101110111011101110111011101110111010101000111011101110111011101000110011101110111011101110111011101110111011001010110011001010101010101010110010101000101010101100101011001100110010101010101010001010110011101110111011101110111011101110111011001010111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101111001100110011001100110011001100110111101110111010111010100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000100001111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000011000100011001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001100100010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100100010000100110011001101000101010101010100010001101000100001110110011101110111100010000100001101000100001100110011001101010110011101100011001100110011001101000110011101100110011001110111011001000100010101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000101011001110111011101110111011101110111011101110111010001000111011101110111011101110111011101110111011101110111010001010111011101110111011001000111011101110111011101110111011101110111011001100101010101100110010101010101010101010110010101100110011001100110011001010101010001000110011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101111001100101110111101110111001011110011011101110110111010100110011001100110011000100010001000100010001000100010001000100010001000100010000111011110001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010000100010001000100011010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010001001000110011001100110011001100110011001101000111100001100011010001000100011101100011001100110011001100110011001100110011010001010011001100110011001100110011010001000011010001010101010000110011010101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010100010001000100010000110011001100110011001100110011001100110011001100110011001100110011001100110010001000100011001100100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001010101010101000100010001010111011101110111011101110111011101110110001101010111011101110111011101110111011101110111011101110111001101010111011101110111011001000111011101110111011101110111011101110111011101100110010101010110010101010100010101110111010101100111011001100110011001100101010101000110011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101111001100110011001100111011001011101110111011101110101010100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000011101111000011110000111100010001000100010001000100010001000100010001000100010001000100010000111011110001000100001110111011101110111011101111000011101111000100010000111100010001000011110001000100010001000100010001000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111010000100010001100110011010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100100001001000110011001100110011001100110011001101000100010101010011001100110011010101000011001100110011001100110011001100110011001101000011001100110011001100110011001100110011001100110011001100110100011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101000100010001000100001100110011001100110011001100110011010000110011001100110011001100110011001100110011001000100011001100100011001100110011001100110011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000101010101010101010001000110011101110111011101110111011101110110001101100111011101110111011101110111011101110111011110000110001101100111011101110111010101010111011101110111011101110111011101110111011101110110011001100110010101010100011101110111010101110111011101100111011001100101010101000110011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001101010101010101010101010101010111011101110101011110111101011101010101010101010101010100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001100110011010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010010001100110011001100110011001100110011001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100001100110100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110010101000100010101000011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010101010101010101010101010101010101010001000100011001110111011101110111011101110101010001110111011101110111011101110111011101110111011110000101010001100111011101110111010001010111011101110111011101110111011101110111011101110110011001110110010101000101011101110111010101110111011101110111011101110101010101010101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110101010101010101010101010101010101010101010101111001011101010101010101010101010100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000011101110111011110001000011101110111100001111000100001111000100010001000100010001000100010001000100010001000100010001000011000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100110010001000110011010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100001100110101011101111000011101110111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010001010101010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110011001000110011001100110011001100110011010001000100010001000100010000110011010001010101010101010101010101010101010101010101010101100111011101110111011101110100010101110111011101110111011101110111011101110111011101110100010101110111011101110111010001100111011101110111011101110111011101110111011101110111011101110110010101000111011101110110010101110111011101110111011101110110010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000110010001000110011001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010010001100110011001100110011001100110011001100110011001101000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011001110101010001010101010101010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000110011001100101011001100101010101010101010101010111011101110111011101100011011001110111011101110111011101110111011101110111011101100011010101110110011001110110010001100111011101110111011101110111011101110111011101110111011101110110010001010111011101110110011001110111011101110111011101110110011001010110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000011101110111011101111000011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000110011001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b000100010010001100110011001100110011001100110011001100110011001100110011001100110011001101000011001100110011010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101011001000100010101010100001101000100011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010100010001000100010000110011010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010000110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000101011001100110011001100110011001010101010101010101011101110111011101010011011101110111011101110111011101110111011101110111011101100011011001110111011001110101010001110111011101110111011101110111011101110111011101110111011101110101010001110111011101110101011101110111011101110111011101110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101000010001000110011001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000010010001100110011001000110011001100110011001100110011001100110011001100110011001101000100001100110011010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110110010101010101010101000011001100110101011001100111011001010100010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100101010101010100010001000100010001000100001100110011001100110011010000110011001100110011001100110011001101000011001100110011001101000100010000110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000011010101110110011101100110011001100110011001010101011001110111011101000100011101110111011101110111011101110111011101110111011101010100011001110111011101110101010001110111011101110111011101110111011101110111011101110111011101110101010101110111011101100101011101110111011101110111011101110111011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000011100110010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000110011001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110011001100110010001000110011001000110011001100110100001100110011001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000011001100110011001100110100001100110011001100110011001101000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001010100010001010101010001000011001100110011001100110100010000110011001100110011001100110011001100110011001100110011010001010101010000110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000100010001000100010001010111011101100110011101110110011001100101010101100111011101000101011101110111011101110111011101110111011101110111011101000100011101110111011101110100010101110111011101110111011101110111011101110111011101110111011101100100011001110111011101100101011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110101010101010101010101010101010100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001111000100010001000100001111000100010001000011110001000100010001000100010001000100010001000011100110010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000110011001101000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110011001000100010001000110011001100100011001100110100010000110011001101000100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110010101010100010101010101010101000011001100110010001100110100010001000011001100110011001100110100010001000011001100110100010101010100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010101010100010101000100010000110101011101110111011101110111011001010111011001010111011001000110011101110111011101110111011101110111011101110111011101000101011101110111011101100100010101110111011101110111011101110111011101110111011101110111011101010101011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100011001000110011001100110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110011001100110010001000100011001100110011001100110011001101000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100101011001100110010100110011001100110011001100110101010001000011001100110011001100110100010000110011001100110101010101010011001100110011001100110011001100110011010000110011001100110011001100110011001100110011010001000100010001000100010101000101010101010100010001000100010101110111011101110111011101100110011001100111010001000111011101110111011101110111011101110111011101110111011000110110011101110111011101100011011001110111011101110111011101110111011101110111011101110111011101010101011101110111011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110100001000110011001100110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100011001100110011001000100011001100110011001100110011001101000011001100110011001100110011001100110100010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110110010000110011001100110011001101000101010001000011001100110011001101000100010000110011001101000101010101000011001100110011001100110011001100110011010000110011001100110100001100110011001100110011001100110011010001000101010101010100010101010100010001000100010001010110011101110111011101100110011001100101001101000111011101110111011101110111011101110111011101110111010101000110011101110111011101100011011101110111011101110111011101110111011101110111011101110111011001000110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100011001100110101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000110011001000100011001100110011001100110011001100110011001100110011001100110011001101000100010001000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101100101010000110011001100110011001100110011001100110011001100110011010001010101010000110011001101010101010001000100010000110011001100110011001100110011010000110011001100110100001100110011001100110011001101000100010001000100010001010101010101010101010101000100010001000101010101100111011101110111010101010100001101010111011101110111011101110111011101110111011101110111010001000111011101110111011101010100011101110111011101110111011101110111011101110111011101110111011001010111011101110111010101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100100011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100011001100100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000110011001100100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101100111011101010100010000110011001100110011001100110100010000110011001100110100010101010101001100110011010001000100010001000100010000110011001100110011001100110011010000110011001100110100010000110011001100110011010001000100010001000100010001010101010101010101010101010100010001000100010101010101011001110111010101100100001101010111011101110111011101110111011101110111011101110111010001010111011101110111011101000100011101110111011101110111011101110111011101110111011101110111010101100111011101110110010101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001100100010001100110011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100110011001100100010001000100010001100110011001100100010001000100010001100110010001100110010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101100111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011001000100001100110011010000110011010001000100010000110011001100110101010101010100001100110100010001000100010001000100010001000011001100110011001100110100010000110011001100110100001100110011001100110011010001000100010001000100010001010101010101010101010001010101010101000100010001010101010101100110011001010100010001100111011101110111011101110111011101110111011101110111001101010111011101110111011101000101011101110111011101110111011101110111011101110111011101110110010101100111011101110110010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000110011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000110011001100110011001100110011001100110011001100110010001100100010001100100010001000110010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111010101000100001100110100010000110011010001010101010000110011001101000101011001010100001101000100010001000100010101000100010001000100010000110011001100110100010000110011001101000100001100110011001100110011010001000100010001000100010001000101010101100110010101010101010101010101010101010101010101000101011001010011010001110111011101110111011101110111011101110111011101110110001101100111011101110111011000110110011101110111011101110111011101110111011101110111011101110110010101110111011101110101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011101111000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001101000100010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110011001100110011001100110011001100110011001100110011001100100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011010001000100010001000101011001110110011001100110011101110110011101100111011101100110011001100111011101110111011101110110010101000011010001000100010000110011010101010100001100110011001101010110010101000100001101000100010001010101010001000101010001000100010000110011001101000100010001000011001101000100001100110011001100110011001101000100010001000101010001000100010101010110011001010101011001010101011001010101010101000101010101000100010101110111011101110111011101110111011101110111011101110101010001100111011101110111010100110110011101110111011101110111011101110111011101100110011101110101010101110111011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100011011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000110011010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110011001100100010001000100011001100110011001100110011001100110010001100110010001000100010001100100011001100110011001000110011001100100010001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001101000100010001000100010101100111011101100110011101110110011101100110011101100110011001100110011101110111011101100101010101000100010001000101010000110011010101100101010000110011010101100110010101000011010001010101010101010101010101010101010001010100010000110011001101000100010001000011001101000100001100110011001100110011001101000101010001000101010101000100010101010110011001100110011001100101011001100110010101010101011001000100011001110111011101110111011101110111011101110111011101110100010101110111011101110111010101000111011101110111011101110111011001100110011001110110011101100101011001100110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110011001100110011001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100011001100110010001100110011001000100011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001101000100010001000100010001000110011101110111011101100110011001100110011101100110011101110110011001110111011101100110010101010100010001000101010000110100010101100101001100110100011001100110010100110011010001010101010101010101010101010100010101010100010000110011001101000100010001000011001101000100001100110100001100110011001101000100010101000101010101010101010001010101011001100110011101110110011001110110011001010101010100110100011101110111011101110111011101110111011101110111011101110100010101110111011101110111010001000111011101110111011101110110011101110111011101110111011101100101011001110111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000011110001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010010110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100100011001100110011001100110011001100110010001000100011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110100011001110110011101100110011001100110011001100110011001110110011001110111011001110110011001100101010101010110010000110100011001010100001100110101011001100101010001000011010101010101010101010101010101010101010101010100010000110011001101000100010101000011001101000100001100110100001100110011001101000100010001000101011001010101010101010101010101100110011001100111011001100110011001100110010100110101011101110111011101110111011101110111011101110111011101100100011001110111011101110110001101010111011101110111011001100111011101110111011101110111011101100101011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011110001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100010001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000110011001100110011001100110011001100110011001100110011001000100010001100110010001000110011001100110011001100110010001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011010001010110011101100110011001100110011001100110011001100110011001100110011001110110011001100110011101100110010101010110010000110100011001010011001101000110011001100101010001000100010101010101010101010101010101100110010101010101010000110011010001000101011001000011001101000011010001000100001100110011010001000100010101010101010101010101010101010101011001100110011001100110011001010110011101110110010000110110011101110111011101110111011101110111011101110111011101100100011001110111011101110101001101100111011101110110011101110111011101110111011101110111011101010110011101110111011001100111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010000111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010010010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100100010001000100010001101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001100110011001100110011001100110011001101000011001100110011001100110010001100110010001000100010001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011010001000101011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110010000110101011001000011001101010111011001010100010001000100010101010101010101010101010101010110010101010101010000110011010001010110011001000011010001000100010001000011001100110011001101000101010101100101010101010110010101100110011101110111011101110111011001010110011101110110010001000110011101110111011101110111011101110111011101110111011101010100011101110110011001100100010001100110011001110111011101110111011101110111011101110111011101010110011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010010001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001000100010001101011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000100010001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110100010001000101011001110110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011001100110010000110100010000110011010001100110011001010100001101000101010101010101010101010101010101010101010101010100001100110011010001010110010101000011010001010101010101000011001100110100001100110101011001100110011001100111011001110111011101110111011101110111011101100110011101110101010001000111011101110111011101110111011101110111011101110111011101000100011001100101010101010100010101100111011101110111011101110111011101110111011101110111011001010111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100111011101110111011101110111011101110111011101110111011110001000011110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001000010001000100010001101000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100011001100110011001100110011001000100010001000110010001000100011001100110011001100110011001100100010001000100011001100110011001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110100011001100110011001100110011001100110011001100110011001100101011101100110011001100110011001100110011001100111011001100110001100110011001100110011011001100110010101000100001101000101010101010101010101010101010101010101010101010100001100110011010001010110011001000010010101010101010000110011001100110100010001000101011001110110011101110111011101110111011101110111011101110111011101100110011001100100001101010111011101110111011101110111011101110111011101110111011001000101011001100110011001010011010101110111011101110111011101110111011101110111011101110111011001010111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110010001000100010001101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001100110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100110011001100110011001100100010001000100010001000110010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100100011001101010110011101100111011001100110011001100110010101010101010001000101011001100110011001100110011001100110011001100110011001100101001100110011001100110100011101100110010001000100001101010110011001100110010101010101010101010101011001010100001100110011010101010110011001000011010101010100010000110100010000110011010001000101011001100110011101110111011101110111011101110111011101110111011101100110011001010011010001100111011101110111011101110111011101110111011101110111011000110110011001100110011001010100011001110111011101110111011101110111011101110111011101110111010101100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001101101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001010010001000100010001100110110100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100110011001100100010001000100010001000100010001000100011001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011010001100111011001100110010101010100010001000100001100110011001100110011010001100110011001100110011001100110011001100110011001100101001100110011001100110110011001010101010000110011010001100110011101100101010101010101010101100101010101000100010000110011010101010110011001000011010101010100010000110100010000110011010001000101011001100110011101110111011101110111011101110111011101110111011001100110011001000011010001110111011101110111011101110111011101110111011101110111010101000110011001100110011001000100011001110111011101110111011101110111011101110111011101110111010101100111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100010001000100010001100110101100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100100010001000100010001000100010001000100010001000100010001100100010001000100011001100110011001100110011001000110011001100110011001100100010001000110011001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110100010101010101010000110011001100110011001100110011001100110011001100100011010101100110011001100110011001100110011001100110011001110101001100110011001101010110010101010100010000110011010101100101010101100101011001010110011001100101010101010100001100110100010101100110011001000011010101010100010001000100010000110100010001000100011001100110011101110111011101110111011101110111011101110111011001010110011001000011010101110111011101110111011101110111011101110111011101110111010001010110011001100110010100110101011101110111011101110111011101110111011101110111011101110110010101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110000111011110001000011101111000011101110111100010000111011101110111011101110111011101110111011101110111100010001000011110000111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000011001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001100110100100010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100011001100110010001000100010001100100010001000110011001000100010001000110010001000100010001100110011001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000110100010001000110011001100110011001100110011001100110011001100100001100110011010101010101010101010100010000110100011001100110010101010110011001010101010101100101010101010100001100110100010101100110011001000011010101010101010001000100010001000100010001000101011001010110011001100111011101110111011101110110011001100110011001010110010100110100011001110111011101110111011101110111011101110111011101110110010001100110011001100110010100110110011101110111011101110111011101110111011101110111011101110110011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001110111100001110111011101110111011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000110100011110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100011001000100010001000100010001000100010001100100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000110011001100110011010001010110011001100110011001100110011001100011001100110100011001010101010101000011001100110101011001100110011001100110011001100110011001100110011001010100001100110101011001100110010100110011010101010100010001000100010001000100010001000100010101100110011001100110011001100110011001100111011001100110010101010110010100110100011001110111011101110111011101110111011101110111011101110110010001100110011001100110010001000110011101110111011101110111011101110111011101110111011101110101011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110000111100010001000100010001000100001111000100010001000011101110111100001110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001100110011011110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100011001100110010001000100011001100100010001000100011001100100010001000100010001100100010001000100011001000100011001100110010001100110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001000100011001100110011001100110011001100110011001100110011001100100010001000100011001100110011010001010110011001100110011001010011001100110100010101010101010000110011001101000110011001100110011001100110011001100110011001100110011001010100010001000101011001100110010100110011010101010101010001000100010001000100010101010100010101100110011001100110011001100111011001100110011001100110011001010101010000110100011001100111011101110111011101110111011101110111011101110101010001100110011001100101001101010111011101110111011101110111011101110111011101110111011101100101011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011110001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001100110011011010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100110011001000110011001100110010001100100011001100100010001000100010001000100010001000100010001100110010001100100010001000100010001000110011001000110011001100110011001100110011001000100010001000100010001000100010001000100010001000100010001000100010001100100010001000100011001100110010001100110011001100110011001100110011001100110011001100110011001000100011001100110011001100110011001100110011010101100101010101010011001100110100010101010101010000110011001101010110011001100110011001100110011001100110011001100110011001010100010001000101011001100110011000110100010101010101010101000100010001000100010101010101011001100110011001100110011001100110011001100110011001100110010101010101010001000101010101100110010101010111011101110111011001100111011101110100010101100101010101100101001101010111011101110111011101110111011101110111011101110111011101100101011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110000111011110001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100001110111011101110111011101111000011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000110010010110001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001100110011001100110011001100110010001000100010001000100010001000100010001000100010001000100010001100110011001100100010001000100010001000110011001100110011001100110011001100110011001100110011001100110010001000100010001000100010001000100010001000100011001100100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001000100011001100110011001100100011001100110011010001010101010101010011001100110100010101010100001100110011010001100110011001100111011101110110011001100110011001100110011001010100001101010110011001100110011000110100010101100110010101000100010001000100010101100110011001100110011001100111011101100110011001100110011101100101010101010100010001000101011001100110011001010101011101110110010101100110011001100100010101100101010101010100001101100111011101110111011101110111011101100111011101110111011101010110011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010000111011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001101000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000110010010010001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001100110011001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001000100010001100110011001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001100110010001000110011001100110011010001000100010101000010001000110100010001010100001100110011010001100110011001110111011101110110011001100110011001100110011001010100010001010110011001100110010100110100011001100110011001000100010001000101011001100110010101100111011101110111011101100110011001100110011001100101010101010100010001000101010101100110011001100110011101100101010101100101010101010100010101010101010101010100010001100111011101110111011101110111011101010110011101110111011101010110011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001100100010001100110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000001100100011001100110011001101111000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001100110011001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100011001100110011001100110011001100110011001100110011001100100011001100100010001000100010001100110010001100110011001100110011010001010100010001000011001101000101010101000011010001000100010001100110011101110111011101110111011101110111011101100110011001010101010001100110011001100110010100110101011001100110011001010101010101000101011001100110011001100111011101110111011101100110011001100110011001100101010101010100010001010101010101010110011001100110011001010101010101010101011001010100010101010101011001010100010101100110011101110111011101110111011101100101011001110111011001010111011101110110010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010000100011001100110010001101111000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000110011001100110011001100100010001100110011001100110011001100110011001100110010001000100010001000100010001000110011001100110011001101000101010000110011001101000101010101000011010001000100010101100110011101110111011101110111011101110111011001100110011001010100010101100110011001100110010000110101011101110110011001100110010101010110011001100110011001100111011001110111011001100110011001100110011001100101010101000100010001010101010101010101011001100110011001010101010101010101010101000100010101010101010101000100010101100101011001110110011001100111011101100101010101100111010101010110011001010101010101010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000010100100011001100110010001001101000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100100011001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100011001100110011001100100010001000100010001100110011001100110011001100110011001100110011001000100010001100110011001100110011001100110011001100110011001000110101010000110100010001000100011001110111011101110111011101110111011101110111011101100110011001010100010101100110011001100110010000110110011101110111011101100110011001100110011001100110011001100110011001010101011001100110011001100101010101010101010101000100010001010101011001100110011001100110011001010101010101100101010101000101010101010101010101000100010101010110011001100110011001100110011101100101010101100110010001010110011001010101010001010101011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010011000100010011001100010001001100010011000100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011000100011001100100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100010001100100010001100100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000101010001000100010001000100010101110110011001110111011101110111011101110111011101100110011001010101011001100110011001100110010001000110011101110111011101110110011001100110011001100110011001100110010101010101010101010101011001100101010101010101010101000100010101010101010101010101011001100110010101010101010101100101010101000101010101010101010001000101010101010110011001100110011001100110011001100110010101100101010001100111011001000100010001000101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111001100100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010001000100010001000100010001000100010001000100110011000100010001000100010001000100010001000100010011000100010001000100010001000100010011000100010001000100010011001100110011001100110011001100110001000100010011001100010011000100110011001100010001000100010011001100010011001100010001001100110001000100010001000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011100110010001100110010001001001000100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001000100010001000100010001000100010001000100010001000100011001100110011001100110010001000100010001100110011001100110011001100110011001000100010001000100010001100110011001000110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100011001100110011001110111011101110110011101110111011101100110010101000101011001010101010101100110010001000111011101110111011101110110011001100110011001100110011001100110011001010101010101010101011001010101010101010101010001000100010101010101010101010101010101100110010101010101010101100101010101010101010101010101010001000101011001100101011001100110011001100110011001100110010101010100010101100101010001000100010001000100010001010110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010001000100010001000100010001000100010001000100010001000001100100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001100110011001100010011001100110011001100110001001100110011001100110011000100010001000100010011000100110011000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001000100010001000100010001000100010001000011100110010001100110010001000110111100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000100010001000100010001100110011001100110011001100100010001000100010001000110011001100110011001100100010001000100010001000100010001000110011001100110011001100110011001100110011001100100010001100110011001100110011001100110011001000100011001100110011001100110011001100100011001101000100010001000100010001000100010101100110011001110111011101110111011101110111011101100110010101000100010101010101010101010101001101000111011101110111011101110110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000101011001100101011001100110011001100110011001010101010001000100010001000100010001000100010001000100010001010101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011000100010001000100010001000100010001000100010001000100010001000100010001000010000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010011001100110011000100010001000100010001001100010001000100010001000100110001001100010011000100010001000100110011001100010011000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110001000100010001000100010011000100110011000100010011000100010011000100010001000100010001000100001000010001100110010001000100110100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100010001000110011001000100011001100110011001100100010001000100010001000100010001000110011001100110011001100100010001000100010001000100010001000100010001100110011001100110011001100110011001000100010001100110011001000100010001000110011001100110011001100100011010001000100001100100011001101000100010101000100010001000100010101100110011001100111011001100110011001100111011001100101010001000101010101010101010101010100001101000110011001100111011101110110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000101010101100110011001100110011001100110011001010101010001000100010000110100010001000100010001000100010001000101011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000011110000111011101100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001001100110001000100110001001100110011000100010001000100110001000100010001000010000100010001000100101100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110001000100110011001100110001000100110001000100010001000100010001000100010001000100010001000100010011001100110001000100010011001100110001001100110011000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010011001100010001000100010001000100001000010001100110010001000100101100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110011001100110010001000100011001100110010001000100010001000100010001000100010001000100010001100110011001100110011001100100010001000100010001100100010001000100010001000100011001100100010001100110011001100110011001100110011001000100010001000100011001100110011001100110100010001000100001000110011010001000101010100110100010001000101011001100110011001100110010101010101010101010110011001100100010001000101010101010101010101010100001101000110011001100110011001100110011001100101010101010101010101010101010101010101010101010101011001010101010101010100010001000101010101010101010101010101010101010101010101010101010101010100010101010101010101010100010001000101010101010101011001100110011001100110011001010100010001000100010001000011001101000100010001000100010101010101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101100111100001110111011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100010001001100110011001100010001000010100100010001000100100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010001000100010011000100110001000100010001000100010001000100010011001100110011001100110011001100010001001100010011001100110001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011000100010001000100001010010001000110010001000100100100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110010001000100010001100100010001000100010001000100010001000100010001000100010001100110011001100110011001000100010001000100010001100110010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110010001100110011001100110100010001000011001000110011010001000101010001000100010001000101011001100110010101010101010101010101010101100110011001010100010001010110010101010101010101010100001101010110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101000100010001000101010101010101010101010101010101010101010101010101010101010100010101010101010101010100010001010101010101010101010101100110011001100110010101010100010001000011010000110011001100110100010001000100010101100110011001100110011101110111011101110111011101110111011101110111011101110111011101100111011101111000011101101000100001110111011001100111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000011101111000011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000010100100010001000100100100010001000100010001000100010001000100010001000100010011000100010001000100010001000100010011001100110011001100010011001100110011001100110001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100001100010001000110011001100100100100010001000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001100110010001000100010001000110011001000100010001000100010001000100010001000100011001100110011001100110011001000100010001100110010001000110011001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100100011001100110100010001000011001100110011010101010100010000110011001101000101010101010101010001010101010101010110011001100110011001000100010001010101010101010101010101010100010001010110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101000100010001000101010101010101010101010101010101010101010101010101010101000100010101010101010101010100010001010101010101010101010101100101010101010101010101010100010000110100010001000100010001000100010001000100010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101100111100010000111011101100111100001110110011101100111100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101100110011101110111011101110111011001100110011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011000100010001000100110001000100010001000100010011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011000100010001000100100100010011000100010011001100010011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100101110011001000110011001100100011011110011000100010001000100010001000100010001000100010001000100010001000,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100011001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001000100011001100110011001000110011001100100010001100100010001000100010001000100010001000110011001100110011001100110011001100110011001100110010001000110011001100110010001100110011010001010100010000110011010001000101010001000101010101010101010101100110011001100110010101000100010101010101010101010101010101010011010001010110011001100110010101100110011001010101010101010101010101010101010101010101010101010101010101010101010001000100010001010101010101010101010101010101010101010101010101010101010101000101010101010101010101010100010001010101010101010101010101100110010101010101010101010100010000110011010001000100010001000100010001000100010101010101010101010110011001110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011001100111100010001000100010001000100010001000100010001000100010001000100010001000100001110110011001100110011101110111011101110110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100010011001100110011000100010001000100010001001100110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011000100010001000100011100010011000100010011001100010011000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100110011001100110011001100110011001100110011001100110011000100110000011001000100010001000100011011010001000100010011000100010001000100110011000100010001000100010001000,
	2400'b001100100010001000110010001000100010001000100010001000100010001000100010001000100010001000100010001000110010001000100011001100110011001100110011001100100010001100110010001100100010001000100010001000100010001000110011001100110011001100110011001000110011001100110011001100110011001100100010001100110011001000110011001100110011001100110010001000100011001100110011001100110011001100110011001100110010001100110011001100110011010001010100010000110011010001000100010001000101010101010101010101100110011001100110010101000100010101010101010101010101010101000011010001010101010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001010101010101010101010101010101010101010101010001010101010101000101010101010101010101000100010101010101010101010101010101100101010101010101010101000100010001000100010001000100010001000100010001000100010001010101010101010101011001110111011101110111011101110111011101110111011101110111011101110110011101100111011101110111011001100110011001100110011101110111011101110111100010001000011101111000011101111000100010001000011101100110011001100110011010000111011101100110011001100110011101111000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100010011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100100010001000100011011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000100010001000100010010110001000100010001000100110011001100010011001100110001001100110011000,
	2400'b001000100010001000100011001000100010001000100010001000100010001000100010001000100011001000100010001000110011001100110010001000110011001100100010001100110010001100110010001100110010001000100010001000100010001000110011001100110011001100110011001000100011001100110010001000110011001100110011001100110011001100110011001100110011001100110010001000100010001000110011001100110011001100110011001100110011001100100011001100100011010001010100001100110011010001000100010001010100010001000101011001100110011001100110010001000100010101010100010101010101010101000011010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001010101010101010101010101010101010101010100010001010101010101010101010101010101010101000100010101010101010101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010101010101010101010101011001110111011101110111011101110111011101110111011101110111011101110110011001100111011101110111011101110110011101110110011101110111011101100111011110001000011101110111011001100111100010001000011101110110011001100110011001100111011101100110011001100110011001110111011101110111100010001000100010001000100010001000100010001000100001110111011101111000100010001000100010001000100010001001100110001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001011100110010001000100010011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110010101001000100010001000100010010010001000100010001000100110011001100110011001100110011000100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000110011001100100011001100110010001100110011001100110010001000110011001100100010001100110011001100110011001100110011001100100010001000100010001000110010001000110011001100110010001100100011001100100010001000110011001100110011001100110011001100110011001100110011001100110011001000100010001000110011001100110011001100110011001100110011001100100011001100100011010001000100001100110011010001000100010001000100010001000101010101010101010101010101010001000101010101010100010101010100010001000011010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010101010101010101010101010101010101010101000100010101010101010101010101010101010101010001000100010101010101010101010101010101010101010101010101010101000100010101010101010001000100010001000100010001000101010101010101010101010101011001110111011001100110011101110111011101110111011101110110011001100110011001100110011001100111011101110110011101110110011101110111011101100110011110000111011101100110011001100111011110001000011101100110011001100110011001100110011101110110011001110110011001110111011101110111100010001000100010001000100010001000100010001000100010000111011101110111011101111000100110001000100110000111100010001000100010001001100001100110011110001000100010001000100010001000100010001000100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100000110010001000100010011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000100010001000100010001101111001100010011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001000100011001100110010001100100010001100110010001000110011001100100010001100110011001100110011001100110011001100110010001000100010001000100010001000100011001100110010001000110011001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110010001000100011001100110011001100110011001100110011001000110011001000110011010001000100001100110011010001000100010001000100010001000100010101010101010101010100010001000100010001000100010001000100010001000011010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010101010101010101010101010101010101010001000101010101010101010101010101010101010101010001000100010101010101010101010101010101010101010101010101010101000100010101010101010101000100010001000100010001000101010101010101010101010110011001110110010101010101011001110111011101110111011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101100110011001111000011101100110011001100111011110001000011101100110011001100110011001100111011101110111011001100110011001110111011101110111011101111000100010001000011101111000100010001000100010000111011101110111011101110111100110011001100001100110011110001000100010011001011101100110011010001001100010011001100001100110011110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100000110010001000100010011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111001100100010001000100010001101101001100010011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001000100011001100100011001100100010001100110010001000110011001100110011001100110011001100110011001100110011001100110010001000100010001000100010001000100011001000100010001100110011001000100010001000110011001100110010001000100010001000100010001000100011001100110011001000100011001000100010001100110011001100110011001100110011001000110011001000110011010001000100001100110100010001000100010001000100010001000101010101010101010101010100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010101000101010001000101010101010100010001010101010101010101010101010101010101010101010001000101010101010101010101010101010101010101010101010101010001000100010001010101010101010100010001000100010001000101010101100110011001010101011001100101010101010101011101110111011101100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001111000011101110111011001110111011110001000100001110111011101100110011001100111100001110111011101100110011001110111011101110111011101110111011110001000011101110111011101111000100010001000011101110111011001101000100110011000011101100110011110000111100110011001011101100110100010011001100110011001011101110110011010011001100110001000100010011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010001000100010010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111001100100010001000100010001001011001100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110010001000100010001000100010001000100011001000100011001100110011001000100010001000110011001100100010001000100010001000100010001000100011001100110011001100100011001000100011001100110011001100110011001100110010001100110011001000110011010001000011001100110011010001000100010001000100010001000101010101010101010101000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010101000100010001000101010101000100010101010101010101010101010101010101010101010101010001000101010101010101010101010101010101010101010101010101010001000100010001010101010101010101010001000100010001000101010101010110010101010101010101100101010101010101011001100101011001100110011001100110011001100110011001100110011001110110011001100110011101110111011101110111011101110110011001100111011101110110011101110111011001110111100001110111011101100110011001100111011101110111011001100110011001110111011101110111011101110111011101110111011101100111011101110111011101110111011101100111011001111000100110000111011101110110011001110111100110011000100001111000100110011001100110011000100001110110011010011001100101110110011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010001000100010010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000001100100010001000100010001001011000100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000100011001100110011001100110010001000100010001000100010001000110011001000100011001100110011001000100010001100110011001100100010001000100010001000100011001100110011001100110011001100110011001100110011001000110011001100110011001100110010001100110010001000110011010001000011001100110011010001000100010001000100010001000100010101010101010101000100010001000101010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010001000101010101010101010101010101010101010101010101010101010001000101010101010101010101010101010001000100010001000101010101100101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101100110011001100110011001110110011101100110011001100110011101100110011001100110011001100111011101110111011001100110011001110110011101110111011001110111011101110111011001100110011101110111011001110111011001110111100010000111011110000111011101110111011001110111100010001000100001110111100110011001100110011000100101110110011010001001011101100110011001111001100110011001100110001000100101110111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010001000100010010010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000010000100010001000100010001001001000100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000110011001000110011001100100010001000100010001000100010001000100010001000110011001100110010001000100010001000110011001100100010001000100010001000110011001100110010001100110011001100110011001100110011001100100011001100110011001100100010001100110010001000110011010000110011001100110011010001000100010001000100010001000100010101010101010001000100010001000101010101000101010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001000101010001000100010001000100010001010101010101010101010101010101010101010101010101010100010001010101010101010101010101010101010101010101010101010100010001000101010101010101010101010101010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001110111011101110111011001100110011001110110011001110110011001100111011101110110011001100110011001100110011101100110011001110111011101100110011101110111011101110111011001110111011110000111011101110111011110001001100110010111100001110110011001111000100001110111011101111001100110011001100101110111100001100110100110011000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100010010010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100100010001000100010001000111000100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000100010001100100010001000100010001000100010001000100010001000110011001100110010001000100010001000110010001000100010001100110010001000110011001100110010001000110011001100110011001100110011001100100011001100110011001100100010001100100010001100110100001100110011001100110100010001000100010001000100010001000100010101010101010001000100010001000100010101010101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001010100010001000100010001000100010101010101010101010101010101010101010101010101010101010100010001010101010101010101010101010101010101010101010101010100010001000101010101010101010101010101010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011101110111011101110111011001100111011101110111011101110111011101110111100110101000011101110111011001111000100110000111011101111001100110011001100001110111011001100110011101100110011001100111100010011001100110011000100010011001100001111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100010001000100010001110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010100100010001000100010001000110111100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001000100011001000100011001000100010001000100010001000100010001100110011001100110010001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100100011001100100010001100110011001100110011001100110100010001000100010001000100010001000100010101010100010001000100010001010101010101000101010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001010101010101000100010001000100010101010101010101010101010101010101010101010101010101000100010001010101010101010101010101010101010101010101010101010100010001010101010101010101010101010100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100111011101110111011101110110011101110111011101110111011101110111011101110111011110000111011101110111011101111000011110001000011110001000100110011001100101110110011001100110011001100110011001100110011110011001100110000111011101111000100010001000100010001000100010011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110010001000100010001110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011000110010001000100010001000100110100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001000100011001000100010001000100010001000100010001100110011001100110010001000100010001000100011001000100010001000100010001000100010001000100011001100100011001100110011001100110011001100110010001000110011001000110011001100100010001100110011001100110011001100110011010001000100010001000100010001000100010101010100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000100010001010101010101000100010001010101010001010101010101010101010001000100010001000100010101000100010101010101010101010101010101010101010101010101010101000100010001010101010101010101010101010100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101100110011001010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111100001110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011110000111011101110111100010001000011001100110011001100111011101111000100010000111011101110111011101110111011110000111011101110111100010001000100001110111011101110111011101111000100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110010001000100010001001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001011100110010001000100010001000100101100110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001100100010001000100011001100110011001100110010001000100010001000100011001000100010001000100010001000100010001000110010001000110011001100110011001100110011001100110010001000100011001000110011001100100011001100110011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001010100010001000100010001010101010101010101010101010101010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101000100010001010101010101010101010101010100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110100010011000011101110110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010000111011101110111011101111000100010001001100110011001100010001001100110011001100110011001100110011001100110011001100101110011001000100010001001111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001000010001000100010001000100100100010011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000110010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100100010001000100010001000100010001000100010001000100010001000110011001100110010001000110011001100110011001100110011001100110010001000100010001000110011001000100011001100110011001100110011001100110100010001000100001100110011001100110011001100100011001100110100010001000100010101010101010101010100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000100010101010101010101010101010101010101010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101000100010101010101010101010101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110000111011101110111100001110111011101111000011101110111011101110111011101110111011101110111011101110111100010000111011101111000100010000111011110001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110000011001000100010001001101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100001010011001100100011001100100011100010011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001100110010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100100010001000100010001000100010001000100010001100100010001000110011001100110011001000110011001100110011001100110011001100110010001000100010001100110011001000100011001100110011001100110011001100110011010000110011001100110011001100110011001000100011001100110011001100110100010001000101010101000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001000101010001000100010101010101010101010101010101010100010001000100010001000100010000110100010101010101010101010101010101010101010101010101010001000100010101010101010101010101010101010100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111100001110111011101111000011101110111011101110111011101110111011101110111100010001000100001110111011101110111100010000111011101110111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110000011001000100010001001011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010011001100110011001100110011011110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001000110011001100110011001100100010001000100010001000100010001000100011001100100010001100110010001000110011001100110011001100110011001100110011001100110010001000100010001100110011001000110011001100110011001100110011001100110100010001000100010001000100010001000011001100110011001100110011001100110011001101000100010001000101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010001000100010001010100010001000101010101010101010101010101010101010100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010001000101010101010101010101010101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000011101111000100010001000011110000111100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001101010000011001000100010001001001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101100011001100110011001100110011011010011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001100100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100010001000110011001100110011001100100010001000100010001000100010001000100011001100110010001000110010001000100011001100110011001100110011001100110011001100110010001000100010001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000011001100110011001101000011001100110011001100110100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000101010101010101010101010101010101010101010101010101010101010100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010001000101010101010101010101010101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101010101010101010101011001010110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001001100110011001100110011001100110011001101010000011001000100010001000111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101110011001100110011001100110011011010011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000110011001100110011001100100010001000100010001000100010001100110011001100110010001000100010001000100010001100110011001100110011001100110011001100110010001000100010001100110011001100110011001101000011001100110011001100110011010001000100010001000100010001000100010001000011001100110011001100110011001100110011001100110011001100110011001100110100010001000101010101010101010101010101010101010101010101010101010101010101010001000100010001000100010001000100010101010101010101010101010101010101010101010100010001000011001100110011001101000100010101010101010101010101010101010101010101010100010001000101010101010101010101010101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101011001010101010101100110010101100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110101010100110011001101010000011001000100010001000111000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000011001100110011001100110011010110011001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001100110011001100110011001100100010001000100010001000110010001000110011001100110011001000100010001000100011001100110011001100110011001100110011001100100010001000100010001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100010001000100001100110100010001000100001100110011010000110011001100110011001000100010001000110101010101010101010101010101010101010101010101010101010101010100010001000011001100110100010001000100010001010101010101010101010101010101010101010100001100110011001100110011001100110100010101010101010101010101010101010101010101010100010001010101010101010101010101010101010101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110010101100110011001100110010101010101011001100101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110000100001000100010001000101000101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001101010011001100110011001100110011001100110011001100110101010100110101010101010101010101010011010101010101010101010101010101010101010101010101001100110011010101010101010100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000110011001100100010010010001001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100011001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001100110011001100110011001100100010001000100010001000110010001000110011001100110011001000110011001000110011001100110011001100110011001100110011001100100010001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000011001100110011001100110100010000110010001100100010001000110100010101010101010101010101010101010100010001000100010001000011001100110011001100110011001100110011010001000100010001010101010101000100010001000011001100110011001100110011001100100011010001000101010101010101010101010101010101010100010001010101010101010101010101010101010101010101010101010101010101010101010101010110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100110011001100110011001100110011001100110011001100110011001110111011101110110011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001000100010001001100110000100001000100010001000100111100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010011001100110011010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101001100110010001000100010001110001001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100011001000110010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100011001100110011001100110011001100100010001000100010001000100010001100110011001100110011001001000101001000110011001100110011001100110011001100110011001000100010001000100011001100110011001100110011001100110010001101000011001100110011001100110011001100110011001100110011001100110011001101000011010001000011010001000010001000110100001100100010001000100010001000100011010001000100010001000100010001000100010001000100010001000100010000110011001100110011001100110011001101000100010001000100010000110011001100110011001100110011001000110011001100110011010001000100010001000101010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010110011001100110011001100101010101010101010101010101011001100110011001100110011001100101010101010101011001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001110111011110001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100010011001100110000100001000100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101001100110011001101010101001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110101010101010011001101010011010100110011001100110011001100110011001100110011001100110011001100110010101001100110010001000100010001101111001100110011001100110011001100110011001100110011001,
	2400'b001000100010001000100010001000100010001000100010001000110011001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000100011001100110011001100110011001100100010001000100010001000100011010000100010001100100011001100100011001100110010001100110011001100110011001100110011001000100010001000100011001100100011001100110011001100110010001000110011001100110011001100110011001100110011001100110100001100110011001100110011010000110011010001000011001000110011001100100010001000100010001100110011001100110011001100110100010001000100010001000100010001000100010000110011001100110011010000110010001000110100001100110100010000110100010001000011001101000011001100110011001000100010001100110100010001000100010001000100010000110011001101000101010101010101010101010100010001000101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111010101111001101010000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000100001000100010001000100110100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111001100110010001000100011001101111010101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001000110011001100110011001100110011001000100010001000100010001000100011001100100010001100100011001100100010001100110011001100110011001100110011001100110011001000100010001000100011001000110011001100110011001100110010001000110011001100110011001100110011001100110011001101000011001100110011001100110011001100110011001100110011001100110011001100100011001000100010001100110011001100110011001100110011010001000100010001010101010101000100010001000100010001000011001101000011001100110100001100110011001101000100010001000011001100110011001101000011001100110011010001000100010001000100010001000100010001000100010001000100010101010100010001000100010001010110011001110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011110000111010101100111011110000111011101110111011101110111011101110111011101100110011001100110011001100110011001100111011101110110011001110111011101101000011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011001100110011001100110011001100110011001100110011001100010001001100110011001100110011000100010001001100110011001100110001001100110001000100110001000100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101001000100010001000100101100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100111001100110010001000100010001101101010101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100010001000100010001000100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110011001100100010001000100010001000100010001100110011001100110011001100110010001100110011001100110011001100110011001100110011001000100010001000100010001100110011001100110011001100110010001000110011001100110011001100110011001100110011010000110011001100110011001100110011001100110100001100110011001100110011001100110011001100110011001100110100010001000100010001000100001101000100010001000100010001000100010001000100010001000100010001000100010101000100010001000100010001000100010001000100010001000100010001010101010001010101010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011001100111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110110011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110001000100110011001100110011001100110011001100110011001100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001100110011001100010001000100010001001100010001001100110011001100110011001100110011001100110011001100110010101001000100010001000100101101010101010100110011010100110011001101010101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000001100110010001000100010001101011010101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000100011001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010001100110011001100110011001100110010001100110010001000100010001000110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100010001000100011001100110011001000110011001100110011001000110011001100110011001100110011001100110100010001000100010001000100001100110100010001000100010000110100010000110011010001000100010000110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111100010000111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011000100010011000100110011001100110011001100110011001100110011001100110001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110001000100010001001100110011001100010011001100110101010101010101010101010101010101010100111001000100010001000100100100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010000110010001000100010001101001001101010101010101010101010101010101010101010101010,
	2400'b001000100010001000100010001000110011001100100011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100001100110011001000100010001100110011001101000100010001000100010101010100010001010100001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010001000100010001000100010001000101010101000100010101000100010000110100010001000100010001000100010101010101010101010101010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010001000101010101000100010001000100010001010101010101010101010101010101010101010100010001000100010001010100010001000100010001000100010101010101010101010110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110001000100010011001100110011001100110011001100110011001100110011001100110101001100110011010101010101010100110011010101010101010101010101010101010101010101010111000001000100010001000100100100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010100110010001000100010001000111000101010101010101010101010101010101010101010101010,
	2400'b001000100010001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011001100110011001101000011010001000100010101010101010101010100001100110100010001000101010100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000101010101000100010001000100010001000100010001000100010001000101010101010100010001000100010001000100010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011110001000100010001000100010001000100010001000100010001000100010001000011101110111011101111000100001110111011101110111011101110111100010001000100010001000100010001000100010001000100110011001100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111001001000100010001000100011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010100110010001000100010001000110111101010101010101010101010101010101010101010101010,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101000100010001000100010001000100001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000100010101000101010101000100010001000100010000110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010001000100010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100001110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001001100110011010101111001100101110111010101010011001100110011001100110011001100110011001100110011001100110101001100110011001100110101001100110101010101010101001100110011001100110011001100110011001100110011001100110011010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010001100100010001000100010100110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011000100010001000100010001000110110101010101010101010101010101010101010101010101010,
	2400'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100010001000100010001000100010001000100010001000100010001000011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011001100110011001100110100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010100010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010100010101010101010001010101010101010110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110101011110111011101110010111010101010011001100110011001100110011001101010101010101010011001100110011001100110011010101010011001100110101010101010101010101010101001100110011001100110101010101010101001100110011001101010011001100110101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001100100010001000100010100010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010011100100010001000100010001000110101101010101010101010101010101010101010101010101010,
	2400'b001100110011001100110011001100110011001100110100010001000011001100110011001100110011001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110011001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001101010101011110111101101110010111011101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101010101010011001100110011001100110011010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010000010001001000100010011110111010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011100110010001100110011001000110100100110011010100110011001101010101010101010101010,
	2400'b001100110011001100110011001101000100001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001100110100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101000100010001000100010001000101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011001100110011001110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011010101010011001100110011001100110011001101010101011110111011101110111001011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010011010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010101010101010101010010100010001001000010010011010111010101110101010101010111011101110101010101010101010101010101010101110101011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100110010001000100010001000110100100010101001100110011001101010101010101010101010,
	2400'b001100110011001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101000100010001000100010001000100010001000100010001000100010001000100010101010101010101000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001110111011101110111011101100111011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010001000100010011001100110011001100110011010101010101010100110011001100110011010101010101011110011011101110111001011101010101010101010101010101010101010101010011001100110101010101010101010101010101010101010101010101010101010101010101010101010101001100010001001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101010111011101010101011011000010001001000010001011010111011101110101010101010111011101010101010101010101011101110101011101010101010101110111011101110101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001000010001000100010001000110100100110111010101010101010101010101010101010101010,
	2400'b001101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101010101010101010101010001000100010001000100010001000100010001010100010101010101010101010101010101000100010001000100010001000100010001000101010101010101010101010101010101000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011101110111011101100111011101100110011001100110011001100110011001100110011001100110011101110111011101100110011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001101010101010100110011001100110011001101010101011110111011101110111001011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010111011101110111011101110111011101010111011011000010001000100010001010110111011101110111011101110101010101110101010101010111011101110111011101010101010101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010101010101010101010101010101011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010011001000100010001000110011100010111011101110111011101110111011101110111011,
	2400'b001100110011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101010101010101010101010101010001010100010001000100010001010101010101000100010001010100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110010101100110011001100110011001100110011001100110011001010101010101010101011001100110011101110111011101110111011101110111011001100110011001100110011001100110011001110111011101110111011001110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100001110111100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011010100110011001100110011001100110101010100110011001100110011001100110101011110111101110110111001011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010111011101110101011101110111011101110111011011100010001000100100001010010101011101110111011101110011001101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100011001000100010001000110011011110111011101110111011101110111011101110111011,
	2400'b001101000011010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101000100010001000100010101010101010001010101010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001010101011001110111011101110111011101110111011101110111011101110111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111100010001000100010001000100010001000100010001000100010001001100110011001100110101001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001101010111011101010011001100110011001100110011001100110101001100110011001101010101100110111101110110111011011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010101010101010101010101010101010101010100110011001100110011010101010011001101010101010011100100001000100100001001110101010101010101010101010001001100110011010100110011010100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101010111010101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101001110011001000100010001000110011011010111011101110111011101110111011101110111011,
	2400'b010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010001010100010001010101010101010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001110110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100110011001100110011001100110011010101110101010100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110101001100110101010101010101100110111101110110111011100101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100001111001100110101010101010101010101010101010101010011001101010101010100110101010100110011010100100100001000100010001001110101011101110111011101110011001101010101010100110101010101010101010100110011001100110011001100110011001100110011010100110011010101010011001101010101010101010101010101010101010101010101010101010101010101110101011101110101011101010101011101110101010101110101011101110101010101010101010101010101010101010101010101010101010101010101010101010111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101010101010101010101010101010101110111011101110111011101110111011101110101010101010111010101010111011101010101010101010101010101010000011001000100011001000100011011010111011101110111011101110111011101110111011,
	2400'b010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010101000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110010101010110010101010110011001100110011001100110011101110111011001100110011001100111011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011010101010101001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011110111101110110111011100101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001001101010101010101010111011101110111010101010101010101010101010101010111011101110111011101000110001000100010001001010011011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110101010101110101011101110111011101010101011101110101010101010101010101010101010101010101010101010101010101010101010101010111011101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101110000011001000110011001000100011010110101011101110111011101110111011101110111011,
	2400'b010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000100010001000100010101010100010001010101010101010101010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010101010101010100010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101100110011001100110011001100110011001100110011001100110011001100111011101110111011001110110011001100110011001100110011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100110011001100110011001100110101010101010101010101110101001100110011001100110101010101010101010100110001000100110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011110111101110110111001100101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101101000001000100010001001010001011101110101011101110111011101110111010101010101010101010101011101010111011101110101010101010111010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101010111011101110101011101110111011101010111011101110101010101010010100001000100011001000100011010110101011101110111011101110111011101110111011,
	2400'b010001000100010001000100010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001000101010101010101010101010101010101010101010001010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101011001100110011001100110011001100110011001100110011101110111011001100111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011101110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101100110111101110110111011100101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101010001000100010001001001111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101011101110111011101110111011101110111011101110111010101010111010101010111010101010101010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101011101110101010101010101010101010100101001000100010001000100011010010011011101110111011101110111011101110111011,
	2400'b010001000100010001000100010001000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001010101010101100110010101010101011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001010101010101010101010101100101010101010101010101010101010101010101010101010110010101010101011001100110011001100110011001100110011001100110011001110111011001100110011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100001110111100010001001100110011010101010101010101010011001100110011001100110011010101010111011101110101010101010101010101010101010101010101010101010101010100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010111100110111101110110111011100101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101100001000100010001000101101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001000100010001000100011010010001011101110111011101110101010101110111011,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001010101010101010101010101010110010101010101010101010101011001100110010101010101010101010101010101010110010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000011101100110011001100110011101111000100010001001100110001000100110101010101010101010101110111011101110111011101110111011101110101010101010101011101110111011101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010111100110111101101110111001011101110101010101010101010101010101010101010101010101010101010101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101110001000100010001000101011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100010011010101110111011101110111011101110111011101110111011101110111011101110111010101010101010101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001100100010001000100011001101111011101010101011101010101011101010101010,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101010110010101010101011001100101010101010101010101010101010101100110010101010101010101010110010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011110001000011101110111011101110111011101110111011101110111011101100110011001100110011001110111011101110111100010001000100010011001101010111011101110111011101110111011101010101010101010101010101010101010101110111011101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101011110111011101110111001011101010101010101010101010101010101010101010101010101010101010101010011000100110001000100010001000100110001001100110011001100110001000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101110010000100010001000101001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010100110001000100010001000100110101011101110111011101110111011101110111010101110101001100110101001100010011001100110101010101010111011101110111011101110111010101010111010101010111011101010111010101110101010101010101011101110101011101010111011101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010100111001100100010001000100011001101111010101010101010101010101010101010101010,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101011001010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000100010000111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010011001100110011001101010101010101010101010101010111011101111001100110011001100101110111011101110111011101110111010101010101010101010101010101010101010101010101010101010101001101010101001101010011001100110011001100110011001100110011001100110011001101010101011110011011101110011001011101010101010101010101010101010101010101010101010101010101010101010011000100110001001101010101001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110000010000100010001000101001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101001100010001000100010001000100010001001101010101010101010011001101010011001100110001000100010001000100010001000100010011001100110101010101010101010101010011000100010011000100010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010101010101011101110101010101010101010101010101000001100100010001000100010001101101010101010101010101010101010101010101010,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010011010101010101010101010111011101110111011101110111011101110111100110011001100110010111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010101010101010101011110011001100101110111011101010101010101010101010101010101010101010101010101010101010101010101001100110011000100110101010101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010010000100010001000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001101010101001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100010001001100010001000100010001000100010001000100010001001100110101010101010011001100110011001100110011001100110011001100110011001100110101011110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110011001101010101010101110111011101110111011101110111010101110101010101010101010101010101001010000100010001000100010001101011011101110111011101110111011101110111011,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001001100110011000100010001000100001111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100110011010101010101010101010101010101010101010101010111011101110111011101110111011101111001100110011001100110011001011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101111001100101110111011101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011000100010001000100111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110101010101010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010001000100001110111011110001000011110000111100001111000100010001000100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001010101110111011101110111011101110111011101110111010101010101010101010101010101010101010100110001000100110011000100110111100101110111011101110111011101110101010101010101010101010101001010000100010001000100010001101001010101110111010101010101011101110111011,
	2400'b011001100110011001100101010101010110011001100110010101100110011001100110011001100110011001100110011001100110011001100101011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100111011101100110011001100110011101100110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001001100110011001100110101010101010101010101010101001100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100110011010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111100110011001100101111001100101110111100110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110010111011101110111010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100000100010001000100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101010101010101001100110001000100010001000100010001000100010001000100010001000100010001000011101110111100010000111100001111000011101110111011101111000011101110111100001110111011101111000100010001000100001110111011110000111011101110111011101110111011110000111011101110111100010001000100010001001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011010101010101010101010101010101010101001010000100010001000100010001101001001101010101010101010101010101010101010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101100110011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011101110111011101110111011101110111011101110110011001110111011101110110011101110111011101110111011101110110011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010011001100110011001100110011010101010101001100110011001100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001001100110101010101010111011101110111011101110111011101110111011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110011001100110011001100110010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100100000100010001000100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110001000100010001000100010001000100010001000100010001000100010001000011110001000100001110111100001110111011101111000011101110111011101110111100010000111011101110111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100110011001101010101001010100100010001000100010001000111000101010101010101010101010101010101010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101011001100110011101100110011001100110011001100110011001100110011001100110011001110111011101110110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010011001101010101010101110111011101110111011101110111011101110111011101110111011101010101011101010111011101110101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100110010111011101110111011110011001100101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100101000100010001000100100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010101001100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101111000100010000111011101110111011101111000011101110111100001111000011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111100010000111011101111000100010000111011101110111011101111000100010001000100010001000010100100010001000100010001000110111101010101010101010101010101010101010,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001110101011001110110011101100110011001100110011001100110011101110111011101110111011101110111011101100111011101110111011101110111011001110111011101100110011101100111011101110111011001110111011101110111011001100110011001110111011101110110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000011110001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010011001101010101010101010101011101110111011101110111011101110111011101010101011101110111011101010101011101110111011101110111011101110111011101110101011101110111011101110111011101110101011101110111100110011001100110011001011101110111011101110111100110010111011101110111011101110101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110000100010001000100100111101010101010101010101010101010101010101010101011101110111011101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000011110001000100010001000100010000111011101110111011101111000100001110111011110000111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010100110010001000100010001000110110100110011001100110011001100110011001,
	2400'b011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110111011101110101011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100110101010101010111011101110111011101110111011101110111011101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010111011101010111011101110111010101010111011110011001100110010111010101110111011101110111100101110101010101110111011101010101010101010101011101110101011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110010110001000010001000100100110101110111010101010101010101010101010101010101010101010101011101110111010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110000111011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000110101100010001000100010001000100010001000,
	2400'b011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101100110011001100110011001110110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111100010001000100010001000100010001000100010001000100010001000100010011001100110011000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101110111011110001000100010001000100010001000100010011001101010101010101110111011101110111011101010101011101110111011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110101010101010101010101010111011101010101010101010101010101010111011101010101010101010101010101010101010101110101011101110111011101111001011101110111100110010111011101110111011101110111011101110111011101110111010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010111001000010001000100010101101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111100010000111011110000111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000110101011101110111011101110111011101111000,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100111011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100010000111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010011001100110011001101010101010101010111010101110111010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101011101110111010101010101010101010111011101010101011101110111011101110101010101010101011101110101010101110111010101110101010101010101011101110111011101110111010101010101011101010111010101010111010101010111011101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111001001000010001000100010100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111100101110111100110010111011101010011001100110011001100110011001100110011001101010101010101010101001100110101001100110101001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000100101011101110111011101110111011110001000,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011000100110011001100110011001100110011000100110001000100010001000100010000111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001001100010001000100010001000100110011001100110101010101010111010101010101010101010101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101010101010101010101010101010101010101010101011101110111010101010101010101110111011101110111011101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111010101010111010101110111011101010101010101110111011101110111011101110111011101110111011101110111011101110111011101110111010001100010001000100010100101010111011101110111011101110111011101110111010101010101010101010101011101110101011101110111011101110101010101010101010101010101010101110111011110011001100110011001100110010111011101110111011101010101010101110111011101110111011101110101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011000100010001000100010001000100010001000011101110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000100100011101110111011101110111011101110111,
	2400'b011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111100010001000100010001000100001110111100001110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001001100010001000100010001000100010001000100010011001100110101010101010101010101010101010101010101001101010011010101010101010101010101010101010101010101010101010101010101001100110011001100110011010101010101010101010101010101010101001100110101010100110101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101010101010101010101010101110101010101010101010101010101010101010101010101010111011101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010001100010001000100010011101010111011101110111011101110111010101010101011101110101010101010101010101010111011101010101011101110101010101010101010101010101010101010101011101111001100110011001100101110111011101110111011101110111010101010101010101110111011110010111011101110111011101110111010101110111011101110111010101010101010101010101010100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010011000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011000110010001000100010001000100100011101111000011101110111011101110111,
	2400'b011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010000111100001110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001111000100001110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101001100110011010100110011001100110011001101010011001100110011010101010011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111010010000010001000100100010100110111011101110111011101110111011101010111011101110101010101010101010101010111011101010101010101110101010101010101010101010101010101110111011101110111011101110111100110010111011101110111011101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101010101011101010101010101010101010101010101001100110011001100110011001100110011010101010011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001001100110011001100110001000100010001000100010001000100010001000100010001000100001110111011101110111011101000010001000100010001000100100011101111000100010001000100010000111,
	2400'b011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101110111011101110101010101110111011101110111011101110111011101110111011101110111011010100100010001000100010100010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101010101011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110101010101010101010101010101010101010101010101010011001100110011001101010111010100110011001100110101001100110011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011101000010001000100010001000100011011110001000100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111100001110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010101010100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101011101010101011101110111011101110111011101110111011101110111011101110111011101010101010101110111011101110111011101010101010010100100010001000100010011110101010101010101010101010101001100110101010101010011001101010101001100110101001100110011010101010101010101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101011101110101010101010111011101110111010101010101001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010111011101010101010101010101001100110011001100110011001100110011001100110011001100110011001101010101010100110011001100110011000100010011000100010001000100010001000100001010010001000100010001000100011011110011001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010000111100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100110011010101010111011101110101001100110011001100110011001100110011001100110011001100110011010110011001011101010101010100110011001101010011001100110101010100110011010101010011001101010101010101010101010100110011010101010101010101010101010101010011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010111011101110111011101110111011101110111011101110111011101110111011101110111011101110101010101010101010011000100010001000100010011010101010101010101001100110011001100110011010101010011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101010101010111011101110111011101110111011101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110101010101010101010101010101001100110011001100110011001100010001000100010001000100001100010001000100010001000100010011110101001101010011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000011101111000100010000111011101110111011101111000100010001000100010001000100110011001100110011001101010011001100110011001100110011001100110011000100010001000011101110111011101110111011101110111011101110111011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100110101010101110111010101010011001100110011001100110011001100110011001100110011010101111001011101010011001100110011001100110011001100110011001100110011001101010101010100110101001101010101001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101011101110111011101110111011101110111011101110111011101110111010101010101010101010101010011100100010001000100010011010011010101010011001100110011001100110011001100110011001100110011001101010011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010100110101010101010101010101010101010100110011001100110011001100110011001100110011001100110011010101010101001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011010101010011001100110011010101010101010101010101010101010101010101010101010101010101011101010101010101010101010100110011001100110011001100110011001100110011000100001100011001000100010001000100010011010011001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001100111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001001100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000011101110111011101110111011101110111011101110111011101110111011110001000100110011001100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110001001100110011010101111001011101010011001100110011001100110011001100110011001100110011001100110011010100110011001100110011010100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011101110111011101110111011101110111011101110111011101010101010101010101010100000110010001000100010010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100101110011001000100010001000100010010110001001100110011001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001001100110011001100110011000100010011000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011001100110011001101010111010100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001101010011001100110011001101010011010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101110111011101110111011101010111011101010101010101010101010100000110010001000100010010010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000011001000100010001000100010010010001000100110001000100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011101110111100010001001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001101010101010100110011001100110011000100010001000100010001000100110011001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000110010001000100010010010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000011001000100010001000100010010010001000100010001001100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011101110110011001100110011101100111011101100111011101100110011001110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100111011110001001101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011000100001110111011101110111011101110111011001110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010001000100010001000100010001000100010011001100110011000100010001000100010001000100010001000100010001000100010001001101110111010100110011001100110001001100010001000100010001000100010001001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100000110001001000100010001110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000100010001000100010001101111000100010001000100110011001,
	2400'b011001100110011001100110011001100110011001110110011001100111011101100110011001100110011001100111011001110111011101110111011101100110011101100110011101110110011001110110011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011110001001100110011001101010101010101010101011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010011000011101110111011110000111011101110111011101100110011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100001111000100010000111011101110111011101110111011101110111011101110111011101110111100010001000011101110111011101110111011101110111011101110111011101110111011110000111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001010110011001011101010011001100110011001100010011001100110011001100110011001100110011001101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010100110011001100110011001100110101001101010101010101010101010101010101010101010101001100110011001100001000010001000100010001110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001001100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000100010001000100010001101111000100010001000100110011001,
	2400'b011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100111011001100110011101110110011001100110011001100110011001110110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100111011001100111011101110111100010000111100010001000011101110111011101110111011101110110011001100110011001100110011001110111100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011000100010000111011101110111011101110111011101100110011001100110011101110111011101110111011101110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110110011101110111011001110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000011110001000011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011010110011011100101110101001100110011001100110011001100110011001100110011001100110011001100110011010101010101001100110011001100110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101000010001000100010001101111001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100001000100010001000100010001101111000100110011001100010011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101100110011001110110011001110110011001100110011001100110011001100101010101010101010101010100010101010101010001010101010001000100010101010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110010101010101011001100111011101110111011101110111011101110111011101111000011101110111011101110111011101110111011001100110011001100110011001110111011110001001100110101010101010101011101110101010101010101010101010101010101010101010101010111011101110101010101010011001100010001000011101110110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101110111100010011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011011110111101101110010111010101010101001100110011001100110101001100110011001100110011001100110011001100110101010101010101010100110011010101010101010101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010001000100010001001101001100110011001100110011001100110011001100110011001100010001001100110011000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110000100001000100010001000100010001001101000100010001000100110011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101110111011101110111011101110111011101110110011101110111011101110111011001100110011001110111011001100110010101010101010001010101010001010101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001010110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001110111100010011001100110011001101010101010101010111011101010111010101010101010101010101010101010101010101010101010101010101010101010101010100110000111011001100110011001100110011001100110011001100110011101110111011101110111011101110111011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000011101110111011101110111011110001000100010001000100010001001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001101010101100110111101110110010111010101010101010101010101010101010101010101010111011101110101010101010101010101010011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101010010001000100010001001101001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010000101001000100010001000100010001001101000100010001000100010011001,
	2400'b011001100110011001100110011001100110011001100110011101100111011101110110011101110111011001110111011101100111011101110111011001110110011101110111011101110111011101110111011101110111011101110111011101100110011001010101010101000100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001110111011101110111011101111000100010000111011110001000100010000111011101110111011101110111011101110111011101110111011101110111100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110000111011101100110011001100110011001100110011001100110011001110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010011001100110011001100110011001100110101100110111101110110010111010101010011001100110011001100110011001101010101010101010101001101010101010101010111011101110111010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001001100110011000100010001001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100101100010001000100010001001101000100110011000100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011001100110011000100010001000100010000101001000100010001000100010001001011000100010001001100110011001,
	2400'b011001100110011001100110011001110110011001110111011101100110011101110111011101110111011101110111011101110111011001110111011101110110011101110111011101110111011101110111011101100110011101110111011101110111011101110111011001100101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001010110011001110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011110001000100110101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110010111011101110110011001100110011001100110011001100110011101110111011101110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001001100110011001100110011001100110011000100010001000100010001000100010001000011101111000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110101100110111101110110010111010100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101010101010011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100010001001100110011000100010001000100010001001100010011001100110011001100101100010001000100010001001011000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110011000100010011001100110001000100010001000100010000101001000100010001000100010001001011000100010001000100110011001,
	2400'b011001100110011001100110011001100110011001110110011101100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001010101011001100111011101110111100010001000100010011001100110011001100110011001100110011001100110001000100010011001100110001000100010011001100110011001101010101001101010101010100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000011101100110011001100110011001100110011001100110011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100001111000100010001000100010001000100010001000100010001000100001110111100010001000011110001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110101100110111101110110010111010100110011001100110011001100110011001100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011000100010001001100010001000100010001000100010011000100010001000100010001000100010001000100010001000100010001000100110011000100010001000100010001001100010001000100101100010001000100010001001011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100010011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100110001000100110001001100010011000100010001000100010000101001000100010001000100010001001010111100010001000100110011001,
	2400'b011001100110011001100110011001100110011001110110011001110110011001110110011001110111011101110110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001010101011001100111011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101001100110011001100110001000100010001000100010001000100010001000100110011001100110011001100010011001100110011001100010000111011101110110011001100111011101100110011001100110011101110111011101110111011101110111011001111000100010001000100001110111011110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110101100110111101110110010111010100110011001100110011001100110011001100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001001100110001000100110001000100010001000100010001000100010000110001000100010001000100010001001000111100010001000100010011001,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001010110011001100110011101110111011101110111100010001000100010001000100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101001100110011001100110011001100010001000100010001001100110011001100110011001100110011001100110011001100110011001100010001000011101110111011101110111011101100110011001100110011101110111011101110111011101110111011001111000100010001000100010000111100010001000100010001000011110000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001101010101100110111101110110010111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110011001100110001000100010011000100010001000100010001001100110001000100110011001100010011001100010001000100010001000100010001000100110011000100110011000100010001000100010001000100010001000100010001000100001110011001000100010001001001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101111000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001001000111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100111011101100110011001100110011001100110011001100111011001110110011001100111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001010101011001100110011101110110011101111000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000011101110111011101110111011101110111011101110111011101110111100001110111100010001000011101111000100010001000100010001000100010001000100010000111100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101010101010101010101100110111101110110110111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001000110111100010001000100010001000100010001000100010001000100010001000100001111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001001000111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110110011001110111011101110111011101100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101010110011001010101011001110111011101100111011101110111100010001000100010011001100110011001100110001000100010001000100010001001100010001000100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011000100010000111011101110111011101110111011101110111100010001001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011110000111100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001101010101100110111101110110110111010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010011001100110011001100110011000100110011001100010001001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001000110111100010001000100010001000100010001000100010001000100001110111011101111000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111011101110111100010001000100010001000100010001000100010001000011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001001000111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101100110011101110111011101110111011101110111011101100111011101100111011101100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001111000100010001000100010011001100001110111011101110111011101110111011110001000100010001000100010001000100110001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011010100110011010101010101001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110101100110111101110110111001011101010101010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110011001000100010001000110110011110000111011110001000100010001000011101110111011101110111011101111000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001001000111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101100110011001100110011001010101010101010101010101010100010001010101010101010101010101010101010101010101010101010101010101010110011001010101010101010100010101111001100010011001100110011010100110101010100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011010101010101010101010111011101110111011101110101011101010111011101010111010101010101011101010101010101010111010101010101010101010101010101010011010101010011010100110011001100110101010101010101010101010011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001101010101100110111101101110110111010101010101010101010011010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110100001000100010001000100110011101110111011101110111011101110111011101110111011101110111011101110111100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011110001000100010000111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000100010001000110111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011001100110011001100101010101010101010101010101010101010101010101010101010101010101010101000101010101010101010101010101010101010110011001100111011101110111100010011001100110101010101010101010100110011001100110011001100010001000100010000111011110001000100010001000100010001000100010001000100010001000100010011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101010101010101010101010101010101001101010101010101010011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111011110001000100010001001100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001101010101100110111011101110010111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010011001100110011001100110011001100110011001100110011001100110001000100010000100001000100010001000100101100001110111011101110111011101110111011101110111011101110111011101110111011101110111011110000111100010001000011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010000111100001110110011001111000011110000111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010000100100010001000110111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001110111011001110111011101100110011101100110011001110110011001100110011001100110011001010101010101010101010101010101010101000101010101010101010101010101010101010101011001010101011001010110011001100110011101111000100010001000100110011001100110101010101010011001100110011001100010001000100001110111011101111000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010100110101010100110101010101010101001100110101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101110101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011110001000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001101010101100110111011101110010111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010011001100110011001100110001000100010010101001000100010001000100101100110011001100110011000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100111011101100110011101100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110110011001100111011101100111011101110111011101110111011101111000011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000110001000100010001000100010001000110111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110110011101110111011101110111011001100110011001100110011001100110011001100110010101010101010101010101010101010101010101010101010101100101010101100110011001100110011001100110011001100110011001110111011110001000100010011001100110011010100110011001100010001000011101110111011101110111100010001000100110011001100110011001100110011001100010001000100010001001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100010001000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001101010101100110111011101110010111010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010100110011010101010101001100110101010100110011001101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100110001000100010001000100010001000100010001000100010000110001000100010000100010101101010101010100110011001100110011001100110011001100110001000011101110111100010001000100010000111011101110111011101110111011101110111011101100110011001110110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011001110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110001000010010001000100010001000110111100010001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011001110111011101110111011001100110011001100110011001100110011001100110011001100110010101010101010101100101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011101110111011110001000100010001000100010001000100010001000100010001000011110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101110111011101110101010101010101010101010101010101010101010101010111011101110111011101110111011101110111010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010111100110111101110110111001011101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110011001100110011001100110011000100010001001100110010110001000100010000100100100100110011001100110011001100110011001100110001001100110001000011110001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100111011001100111011001100110011001100110011001100110011001110111011001100111011101110111011101110111011001110111011101110110011101110111011101100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110110001000010010001000100010001000110110100010000111100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110110011101110111011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101011001100110011001100110011001100101010101010101010101010101011001100110011001100111011101110111011110001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110001000100110011001100110011001100110011001100110011001100110011010101010011001100110101010101010101010101010101010101010101010101010101010101010111010101010101011101010101011101110111011101110111010101010111011101010101010101010111011101110111011101110111011101110111010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100110001000100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010111100110111101110110111001011101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110010111001000100010001000100100100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011001100111011101100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011101100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010000111011101110111011101110111011101110110001000010010001000100010001000110110011101110111100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101100110011001100110011001110111011101110111011101110110011001100110011001100110011001100110011001100110011001100101010001010101010101010101010101010101010101010101010101100110011001100110010101010101010101010101010101010101011001100110011101110111011110001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001100110101001100110101010101010101010101010101010101010101010101010101010101010101011101110101010101010101010101010101010101010101010101010101010101110111011101110101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101010100110011010101010011001100110011001100110011001100110011001100110011010101010101010101010011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011010101010101010101010111100110111101110110110111010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110101000001000100010001000100011100010011001100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100111011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110110011101100110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000100010001000100010001000100110011101110111011110001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110010101010101010101010101010101010101010101000101010101010101010101010101010101100110011001100101011001010101010101010101011001100110011001100110011101110111011101111000100010001000100010001000100010001000100010001000100010011001100110011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110101010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101001100110011001101010101010101010101010101010101010101010101001100110011010101010101010101010101010101010101010101010101010101010101010100110001000100010001000011110001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001101010101010101010101010101010111100111011101110110111001010101010101010101010101010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001101010011001100110011001100110011001100110010111001000100010001000100011011110001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110001000100010001000100010001000100110011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101100110011101110111011101110110011001100110011001100110011001100110011001100110010101010101010101000101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100111011101110111011110001000100010001000100010001000100010001000100010001000100110011001101010101010101010101010101010101010101010011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101100111011111110110111001011101010101010101010011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101001100110011001100110011001101010101001101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011000001100100010000100100010011110011000100010001000100010001001100110011001100110011001100110101001100110011001100010001000100010001000100010001000011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111100001110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110101001000100010001000100010001000100110011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011001100110011101110110011101110110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001110111011101110111011110001000011101111000100010001000100010001000100010001000100110011001100110011010101010101011101010101010101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010011001101010101010101010101010101010101010101010011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110001001100110011001100110011001100110011001100110011010101010101001100110101010101010101010101010101010101010101010101010111100111011111110110111001011101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101001100110101010101010101010101010101010101010101010101010101010100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001001100100010000100100010011110101001100110011001101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011101110111011101110111011101110111011101110111011101110111011101110111100010000111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110100001000100010001000100010001000100110011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101100110011101110111011001100110011101110111011001100110011001100101010101010101010101010101010101010101010101010100010001000101010101010101010101010110011001100110011001100110011001100111011001110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000100110011010101010101011101110111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001101010101010101010101010101010101010101010101010101010101011101010011001101010101010101010101010101010101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010111011101110111100111011101110110111001011101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010000100010000100100010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100010001000100010001000100010001000100001111000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101111000011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110101001000100010001000100010001000100101011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110111011101100110011001100111011101110111011101110111011101110111011001100110011001100110010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001110111011101110111011101110111011101110111011101110111011110001000100010001000100010001000100010011001101010101010101110111011110011001100101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110101010101010101010101010101001101010101010101010101011101010011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110101010100110101010101010101010101010101010101010101010101010101010101010101011101110111011101110111101111011111110110111001011101010101010100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011010101010101010101010101001100110101010101010011001100110011001100110011001100110011001101010101010101010101001100110011001101010101010101010101010101010101010101010101010101010101001101010101010101010101001101010101010010100100010000100100010010110011001101010101010101010101010101010101010101010101010101010101010101010011001100110101010101010101010101010101010101010101001101010011000100010001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110110011101110101001000100010001000100010001000100101011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101100110011001100110011101110110011101110111011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001110110011001100110011001100111011101110111011101110111011101111000100010001000100010001000100010001001100110011010101110111100110011001100110011001100110010111011101110111010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110101010101010101010100110101010101010101010101110011001100110101010101010101010101010101010101010011010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111100111011111110111011001011101010101010101010101001101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001101010101010101010101010101010011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001010100100010000100100010010110101001101010011001101010011001100110011001100110011001100110011001100110011000100010011001100110011001101010011010101010101010101010101010100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011001100110011001100101001000100010001000100010001000100101011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001110111011101110111011101110111011101110110011001100110011001100111011101110111011101110111011001100110011001010101010101010101010101010101010101000101010101000101010101010101010101010110011001100110011001100110011001110111011101110111011101110111011101110111011110001000100010001000100010001000100110011010101110111100110011001100110011001100110111001101110011001100101110111011101110101010101010101001100110011001100110011001100110011001100110011001100110011010100110011010100110011001101010011001101010101010100110011001100110011010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101011101110101010101010101010101010101010101010111100110111101110111011001011101010101010101010101010101010101010101010011010101010101010101010101001101010011001100110101010101010101001100110011001100110011001100110101010101010101010101010101001101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011100100010001000100010010110101010101010101010100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001101010101001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011110001000100010001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011001100110011001100100001000100010001000100010001000100100011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001100110011001100111011001100110011001110110011001100110011101100111011101110111011101110111011101110110011101110111011101110111011101100110011001100110011001010101010001010101010101000100010001000101010101000101010101010110011001100110011001100110011001100111011101110111011101110111011101110111011101110111100010001000100010011001100110101010101010111011101111001100110011001100110011001101110111011101110111011100110011001100101110111010100110011001100110011001100110011001100110011001100110011010100110011001100110011010101010101010100110011010100110011010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111010101010101010101010101010101110111100110111101101110111001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011010011100100001000100010001010110101010101010101010101010011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001001100110011010101010101010101010101010101010101001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110101001000100010001000100010001000100100011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101100111011101110111011101110111011101110111011101110111011101110111011101110110011001100101010101010101010101000100010001010101010101000101011101100101011001010101010101100110011001110110011001110110011101110111011101110111011101110111011101111000100010001001100110101010101010101010101010101011101110111011110011001100110011001100110011011101110111011101110011001100110011001011101110111010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101010100110011001101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110111011101010101010101110111101111011101101110111001011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101010101010101001101010101010100110011010101010101001101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010011010100000100010001000100010010010101010101010101001101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001001100110011001100110101010101010101010101010101010101010101000100010001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111100001110111011101110111011101100111011101110111011001100110011101100100001000100010001000100010001000100100011101110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100110011001110110011101100111011101110111011101110111011101110111011101100110011001110111011101110110011001100110011001100101010101010101010101010101010101010101011110000110010101100110011001100110011001100110011001100110011101110111011101110111011101110111011101111000100010001000100010011001100110011010101010101010101010101010101010101010101010111011101111001100110011001100110011011101110111011101110111001100110011001100110011001100110011001100110011011101110011001100101110111010100110011010100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101010101010101010101010101010101110111100110111011101110010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010011010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110101010101010011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010100000100010001000010010001110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110011000100010001001100110011001100110011001100110011001100110011001100010011001100110011000100010001000100010011001100110011001100110011001100110011001100110001000100010001000011101110111011101110111011101110111011101110111011101111000100010001000100001110111011101111000100010001000100001110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100100001000100010001000100010001000100100011001110111011101110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110110011101110111011001110110011001100110011101110111011101100110011001100110011001100110011001100111011101100110011001110111011101110111011001100110011001100110011001100110011001100110011001100110011001110110011001100111011001100110011001110110011101110111011101110111011001100111011101110111011101110111011101100110011001100110010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011110001000100010011001100110011010101010101010101010101010100110011001100110101010101010101010101110111011101110111011110011001100110010111011101110111011101110111011101110111100110011001101110111011100101110101010100110011001101010101010101010101010101010101010100110011001100110101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011110011001011101110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100000110001001000010001001110001010100110101010101010011001100110011001101010101001100110011001100110011001100110011010100110011010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010100110011001100110001000100001110111011110001000100010011001100110011001100110011001100010000111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101100110011001100110011001100110010101100110010101010101011001100110011001100110011001100110011001100110011001100110011001100100001000100010001000100010001000100100011001110110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100110011001110111011101110111011101110111011001100110011001100111011101110111011001100110011001100110011101100110011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100101010101010101010101010101010101100110011001100110011001010101010101010110011001100110011001100110011001100110011001110111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001101010011001100110011001100110101010101010101010101010101010101010101010101010101010101110111011110011001011101010101010100110011001100110011001100110011001100110011001100110101010101010101001101010101001100110011010101010101010101010101010101010101010101010101010101010101010101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010111011110011001100101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100100110010001000010010001110001010101010101010101010101010101010101010101010101001100110011001100110101010101010101010101010101010101010101010101010101010101010011001100110011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010011001101010101001100110011001100110011001100110011001100110011001100010000111011101110110011001100110011001100110011001110111011101111000100010000111011101110111011101110111011101110111011101110111011101100110011001110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100101010101100110011001100110011001100110011001100110011001100100001000100010001000100010001000100100011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001100111011001100110011001100110011001100110011001100110011001110110011101100110011001110110011101110111011001110111011001110111011101110111011101110111011001100110011101100110011001100110011101100110011001100110011001100110011101100110011101100111011101100111011101100111011001110111011101110111011101110111011101110111011101110111011101110111011101110110011001010101010101010101010101010101010101100110010101010101010101010110010101010110011001100110011001100110011001100110011001110111011101110111100010001000100010001000100010011001100110011001100110011010100110101010100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101011101110111011101110111010101010101010101010011001100110011010100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011010101010011010101010101010101010101010101010101010101010101010101010101011101111001100101110111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010100110011001100110011001100110011001100110011010100101000001001000010010001010001010101010101010101010101010101010101010101010101010101010011001100110101010100110011001100110011010101010101010101010101010101010101010100110011010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100001110111011101110111011101110111011101110111011101110110011001100110011001100111011101110111011110001000100001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000100010001000100010001000100100011001100110011001100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011001110111011101110111011101110111011001110111011101110111011101110110011101100110011001100111011001100110011001100111011101110111011101110111011101110111011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110010101010101011001010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011110001000100010001000100010001000100110011001100110011010101010101010101010011001100110011001100110011000100010001000100010001001100110011001100110011001101010101010101010111011101111001100110010111011101110111010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011010101010011001100110011001100110011010101010101010101010011001101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001000001000100010010001010001011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010011001100110011010101010101010101010101010100110011001101010101010100110011001100110011001100010001000100010001000100010001000100010001000100010001000100001110111100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100101001000100010001000100010001000100011011001100110011101100110,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001110111011001110111011101110110011101110111011101110111011101110110011001100110011001110111011101110111011101110111011101110111011101110110011001110111011101100111011101110111011101110111011101110111011101110111011101110111011001100110011001100110010101010101010101010101010101010101011001010101010101010101010101010101010101100110011001110111011001110111011101110111011101110111011110001000100010001000100010011001100110011010101010011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010011001100110101011101110111011101110111011101110111011101110111011101010101010101010011001101010101010101010101010101010101010101010101010101010101010100110011010101010101010101010101001100110011001100110011001100110011010101010101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001010010001000010010001001111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010100110101010101010101010101010101010101010101001100110011001101010101010101010101001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100010001001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000111011101110111011101110111011101110110011001100110011001100110011001100110011001100111011101110101001000100010001000100010001000100011011110000111100001110111,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001100111011101110111011001100110011001100110011001100110011101110110011101110110011001110111011101100111011101110111011101100111011101110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010110011001100110011001100110011001110111011101110111011101110111100010001000100010001000100010001001100110001000100010001000100010001001100110011001100110011001100110011000100010001000100010001000100010001000100110011001101010101011101110111011101111001100110010111011101110111010101010101010101010101010101010101010100110101010100110011001101010101001100110101010100110011001100110011001100110011001100110011001100110011001100110101010101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101100010001000100010001001101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010011001100110101010101010101010101010101001100110101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001001100110001000100010001000100010001000100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101100110011101100110011101110111011001110111011101100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100101010101010101010101010101010101100110010101010110011001100110011001100110011101110111011110001000100010001000100010001000100010001000100010001000100010001000100010011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001001100110011010101010101010101010101011101110111010101010101010101010101010101010101010100110011010101010011010100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100010001000100010001001101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011101110110011001100110011001100110011001100111011001100110011101100110011101110111011101110111011101110111011101110110011101110111011101110111011001110111011001110110011001110111011101110111011101110111011101110111011101110111011101110111011101100111011101100110011001110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001010101010101100110011001100110011001100110011001100110011001100110011101110111011101110111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000011110001000100010001000100010001000100010011001100110011001100110011001100110101010101010011010100110101001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100010001000100010001001011010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110101010101010101001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010000111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100001001000100010001000100011011110001000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101110111011101110110011001110110011001100110011001100110011001100111011001100111011001110110011001100110011001100110011001100110011001110110011101110111011101110111011101110111011101110111011001110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011110001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001110010001000010010001001001010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100001110111011101110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110110011101110110011001100110011001100110011001100110011001100110011001110110011001100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011110001001100110011001100110011000100010001000100010001000100110011001101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101010101010101010101010101010101010101010101010101010101001110010001000100001001000111001101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110101010101010101010100110011001100110011001100110101010100110101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100110011001110110011001100110011001100110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101111000100110011001100110011001100010001000100110011000100110011001100110011001100110011001101010011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101110101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110000010001000010010001000111001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110101010101010011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001001100110011001100110011001100110011000100010001000100010001000100010001000100110001000100010001000100010001000100001110111011110001000100010001000011101110111100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011101100110011001110110011001100110011101110111011001100110011001110111011101110111011101110111011101110111011101110111011101100111011101110111011101110111011101110111011001110111011101110110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011101110111011101110111011001100110011001100110011001100110011001100110011001100111011101110111011110001001100110011001100110011001100010001000100010011001100110101010100110101010101010101001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011001101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111011101010101010101010101010101010101010101010101010101010101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000010001000010001000100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110101001100110011001100110011001100110011001100110011001100110011010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010110011001100110011001100110011001100110010101100101010101010101010101010101010101010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011001100110011001100110011001110111011001100110011001110111011001100111011001110111011001110111011101110111011101110111011101110111011101110111011101110111011101110111011101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110111011110001001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010101001100110011001100110011001100110011010100110101010101010101010101010101010100110101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010000010000100010001000100101000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100110011010101010101010100110011000100010001000100010001000100010001000100010001000100010001000100010001000100110011001100110001001100010011001100110011001100110011001100110011001100110011001100110001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010101010101010101010101010101011001100110010101010100001100110011010001010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101110110011101100111011101110111011101110110011101110111011101100110011101110110011101110111011101110111011101110111011101110111011101110111011101110111011101110111011001100110011101110110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011110001000100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101001101010101010101010101001101010101010101010101010100110101010101010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010010011000100010001001000100111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101110101010101010101011101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010101010101010101010101010101010101010101010101000011001100110011010001010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011001110111011101110111011101110111011101110110011101100111011101100110011001110110011001100110011001110110011001100111011101110110011001100111011001100111011101110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111100010011001100110011001100110011001100110011001100110011010101010101010101010101001101010101010101010101010101010101010100110011001101010011001100110011001100110011001100110011010100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011010100110011010101010011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101001100110011010101010101010101010101010101010101001100110011010101010101010100110011010101010101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011010101010101010101010011001101010101010101010101010101010101010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010010011000100100010001000100110101010101010101010101010101010111010101010101011101010111011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010111011101110111011101110111011101010101010101010101010101010101010100110011001100110011000100010001000100010001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010011001100010001000100010001000100110001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010101010101010101010101010101010101010100010001000100010001000101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011001110110011101110111011101110110011101100110011101100111011101100111011101110110011001100110011001100110011001100111011001100110011001100111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011101110111011110001000100010001000100010011001100110011001101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110101010101010101010100110011001100110011001100110011001100110011001100110011001100110011010101010011001101010101010101010101010101010111011101110111011101010101010101010101010101010101010100110011001100110011001100110011010101010101001100110101010101010101010101010101010101010101010101010101010100110101010101010101010101010101010100110101001100110011001100110101010101010011001100110011001100110011001101010101010101010101010101010011010101010101010101010101010101010101010100110101010101010101010101010101010101010100100000100100010001000100101101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010101010101010101011001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100101011001010101010101010101010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011110001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010011001101010101010101010101010101010101010101010101011101110111011101110101010101010101010101010011001100110011001100110011001100110011001100110101010100110101001101010101010101010101010101010101010100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110101010101010101001100110011001101010101010100110011001101010101010101010101010101010011001100110101010101010011010101010101010101010100100000100100010001000100101101010101010101010101010101010101010101010101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b010101010101010101010110010101100110011001100110011001100110011001100101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001010101010101010101010101010101010101010101010101010101010101010101011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100111011101100110011101100111011101110111011101110111011101110111011110001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011001100110011001100110101010100110101010100110101001100110011001101010101010101010011001100110101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010011001100110101010100110011001100110011001100110011001100110011001100110011010101010011001100110011001100110011001100110010100000100100010001000100101101010101001101010101010101010011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010101010101001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010101110111011101010101010101010101001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110001000100010001001100010000101001000100010001000100010001000100011011110001000100010001000,
	2400'b011001100110010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110010101010101010101010101010101010110011001010110010101100110011001100110011001100110011001010101010101010101010101010101010101010101010101010110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111011001110111011101110111011101110111011101110111100010001000100010001000100010001000100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101001100110011010101010101010101010011010100110011010101010011001100110101001100110011001101010011001101010101010101010101010101010011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001101010011010101010101011101110111011101010101010100110011001100110011001100110011001100110101010101010101010100110011001100110101001100110100101001000100010001000100100100110011001100110101001100110011001100110011001100110011001100110011001100110011001100110011001101010101011101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110001000100010001000100010001000100010001000100010001001100110101010101010011001100110011001100110011001100110011001100110101010101010101010101010011001100110011001100110011001100110011001100110011001100110010101001000100010001000100010001000100011011110001000100010001000,
	2400'b011001100110011001100110010101010101010101010101010101100110011001100110011001100110011001100110011001100110011001100110011001100101010101010110011001100110011001100110011001100110011001100110011001100101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110111011101110111011101110111011101110111011101110111011101110111100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101110101010101010111011101110101010100110011001100110011001100110011001100110011001100110101001100110011001100110011001100110100110001000100010001000100011100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010100110101001100110101010101010101010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110010101001000100010001000100010001000100011011110001000100010001000,
	2400'b011001100110011001100110011001100101010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101010101010101100110011001100110011001100110011001100110011001100101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001110110011001110111011101110111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110101010100110101001100110101010100110101001101010101001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011010101010101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110101011101110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100110001000100010001000100011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011001100110101010101010101011101110101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001101010011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101010101010100110011001100110000100001000100001001000100010001000100011011110011000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101100111011101110111011101110111011101110111011101111000100010001000100010001000100010001000100010001000100010001000100010001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010011010101010101010100110011001101010101010101010101010100110101001100110011001101010101010101010101010101010101001100110101010101010101010101010101010101010101010101010011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110100110001000100010001000100011100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010101010101010101010101010101010101010101010101010101010101010101010101010011001101010011001100110011001100110011001100110011010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010101010101010101010101010011001100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101001100110011001100110010100001000100001000100100010001000100011011110011000100010001000,
	2400'b011001100110011001100110011001100110011001100110011001010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010101010101100101010101010101010101010110010101010110011001100110011001100110011001100110011001100110011101110111011101110111011101110111011110001000100010001000100010001000100010001000100110011001100110011000100010001000100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001100110011001100110101001100110011010100110011001101010101010101010101001100110011001100110011001100110011010100110101010100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010111001000100010001000100010011110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101001100110011010100110101010100110011001100110011001100110011001100110011001100110011001100110011010101010011001101010011001100110011001100110101010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001100110011001100110010100001000100001001000100010001000100011011110011001100010001000,
	2400'b011001100110011001100110011001100110010101010101010101010101011001100110011001100110010101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001010110011001010101010101010101010101010101010101100101010101010110011001100110011001100110011001100111011101110111011101111000100010001000100010001000100010001000100110011001100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110101010101010011001101010101001100110011010100110011010100110011001100110011001100110011010101010101010101010101010101010101010101010011001101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000100010001000100010011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010101010101010101010011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010101010101010101010101010100110011001101010101001100110011001100110101010100110011010100110101010100110011001100110011001101010101010100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110010100001000100010001000100010001000100011011110011001100110001000,
	2400'b010101010110011001100110010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010101010110011001100110011001100110011001100110011001110111011101110111100010001000100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101001101010101001100110011001100110011001100110011001100110011001100110011010101010101010100110011010101010101001100110011001100110101010101010011001100110011001100110011001100110101010101010101001100110101010101010101010101010101010101010101010101010101010101010011001101010011010101010011001100110011001100110011001100110011000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000100010001000100010011010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110010100000100010001000100010001001000100011011110011001100110001000,
	2400'b010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111100010001000100010001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110101010100110011001101010011001101010101001101010101001100110011010101010011001100110101010101010101001100110011001100110011010101010011010101010101010100110011001100110011001100110011001100110011001100110011001100110101001100110011001100110101010101010101010101010101010101010101010101010101010101010011001100110011001100110011001100110011001100110011001100110001000100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110010110001000100010001000100010010110001000100010001000100010001000100010011001100110011001100110011001100110011001100110011001100110011001100110011001100110011010100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010011001100110011001100110000100000100010001000100010010001000100011100010011001100110011001,
	2400'b010101010101010101010110010101100110011001100110011001100110010101010101010101010101010101010101010101010101010101010110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011101110111100010001001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010101010101010101010101010101010101010101010101010101010101010011001100110101010100110101010100110011001100110011010101010011001100110011001101010011001100110011001100110011010101010101010101010101010101010101010101010101010101010101010100110011001100110011001100110011000100010001001100110001000100010001001100110001000100110011000100010011001100010001001100110011001100110001001100110011000100110011001100110011001100110001000100010001000100010001000100010010110001000100010001000100010010110001000100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101010011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100110011010101010011010101010101010101010101001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000100000100010001000100010001001000100011100010011000100010011000,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		// r_data = r_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		// g_data = g_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		// b_data = b_picture[(y_cnt - y_pin)/5][((x_cnt - x_pin)/5)<<3 +: 8];
		r_data = {{picture[(y_cnt - y_pin)][((x_cnt - x_pin)<<2 +: 4)]}, {4'b0}};
		g_data = {{picture[(y_cnt - y_pin) + Y_WIDTH][((x_cnt - x_pin)<<2 +: 4)]}, {4'b0}};
		b_data = {{picture[(y_cnt - y_pin) + (Y_WIDTH << 1)][((x_cnt - x_pin)<<2 +: 4)]}, {4'b0}};
		// r_data = 8'b0;
		// g_data = 8'b0;
		// b_data = 8'b0;
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule