module red_reverse(
	input [9:0] x_cnt,
	input [9:0] y_cnt,
	input [9:0] x_pin,
	input [9:0] y_pin,
	output [7:0] r_data,
	output [7:0] g_data,
	output [7:0] b_data
);
localparam X_WIDTH = 30;
localparam Y_WIDTH = 50;
localparam [0:149][239:0] picture = {
	240'b111011111111001011101010110000011011000110110011101100111011001010110010101100101011001010110011101100111011001110110011101100111011001110110010101100101011001010110010101100111011001110110011101100111011000110111110111001001111000111101111,
	240'b111100101101111010111101110111111111100011111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100011011101101110001101111011110010,
	240'b111001101011100111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001011100111101000,
	240'b101100111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010110010,
	240'b101000111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110100001,
	240'b101100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101,
	240'b101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011,
	240'b101001011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110100100,
	240'b101011011110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001010101100,
	240'b111000001011101111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001011101011100010,
	240'b111100101101010011000000111011111111111011111110111111011111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111101111111101111111111101110101111001101010111110010,
	240'b111110011111110011011101100111001001101010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001100110100001111000111111110011111001,
	240'b111011111111001111101010110000011011000110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011000110111111111001001111001011101111,
	240'b111100101101111010111101110111111111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111100111011101101110001101111011110001,
	240'b111001101011100111110010111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111100001011100111101000,
	240'b101100111101111011111111111001111001100101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011110010111100101111100011111011001101111101001111111111101110010110010,
	240'b101000111111101011111001100001000100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001010111100100111001110101100110010011110100110110000111111110101111101010100001,
	240'b101100101111111111011111010110110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100001111010111111111010000110010011110101001101011110111000101111111110110001,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100001110010111111110011100101011100010100111101011100110110101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111100100011100001011111111110110110110011101011010110110101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101110011011101001011000111111111111011100001011001110110101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101111111111111000101110100111101001101011100110110101111111110110101,
	240'b101101101111111111010111010110100101010001010010010100000101001001010010010100000101000001010001010100110101010101010101010101010101010101010101010101010101010101010011011010001101101111111111110000111001001001011111110110101111111110110101,
	240'b101101011111111111010111010110100101000001101001100110101011000010101111101001111001010001111010011000000101001101010001010101000101010101010101010101010101010101010101010100010111001011100100111110101100001101101010110110001111111110110101,
	240'b101101011111111111010111010101111000011111100101111111111111111111111111111111111111111111110111111000011011100010000001010110000101000101010100010101010101010101010101010101010100111110000101111111111110110001101100110110001111111110110101,
	240'b101101011111111111010011011111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011001000000101010100010100100101010101010101010101010101001101101000101000001001010101100011110110011111111110110101,
	240'b101101011111111111010111110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111001011001010101000101010101010101010101010101010100010100010101000001011100110110101111111110110101,
	240'b101101011111111111100111111100111111111111111111111111111111111111111111111111111111101111111010111110101111100111111000111111111111111111111111110111010111100001010001010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111110000111110101111111111111111111111111111111111111111111110011001010101111100011111110111111010111001111111101111111111111111111111111110101110000011010100000101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111110000111110101111111111111111111111111111111111111111111101110111000001001101010011110110001011100100111111111111111111111111111111111111111111101110011111110101000001010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111101101111110011111111111111111111111111111111111111111111101110111001101010001010101010101010010011011111110111111111111111111111111111111111111111111111001100110111101010001010101010101010001011100110110101111111110110101,
	240'b101101101111111111101001111101101111111111111111111111111111111111111111111101110111000101001101010101000101010001010011101010001111111011111111111111111111111111111111111111111100111101011100010100110101010001011100110110101111111110110101,
	240'b101101101111111111100001111001111111111111111111111111111111111111111111111101011000011110010001010101110101010001010011010101111011100011111111111111111111111111111111111111111111111110100101010100010101001101011100110110101111111110110101,
	240'b101101101111111111011000110100101111111111111111111111111111111111111111111110011101110111101010100111110101001001010101010100110101101111000110111111111111111111111111111111111111111111110000011100100101000001011100110110101111111110110101,
	240'b101101011111111111010010101100101111111111111111111111111111111111111111111111111101100101110110110101001001010001010000010101010101001001100010110100111111111111111111111111111111111111111111101111000101001001011100110110101111111110110101,
	240'b101101011111111111010010100011001111110111111111111111111111111111111111111111111010110101001010011101101101100110000110010100000101010101010000011100101110111011111111111111111111111111111111111100110111000001011001110110101111111110110101,
	240'b101101011111111111010101011010001110011011111111111111111111111111111111111111111010000101001111010100001000001011011010011110100101000001010101010100011011111011111111111111111111111111111111111111111010101001011000110110101111111110110101,
	240'b101101011111111111010110010101111011011111111111111111111111111111111111111111111011010001010000010101010101000010010000110110000110111101010001010100001010011011111111111111111111111111111111111111111101110101100101110110011111111110110101,
	240'b101101011111111111010111010101100111101111111001111111111111111111111111111111111110010001100101010100010101010101010001100111101101001101100101010011001010110111111111111111111111111111111111111111111111100110000101110101101111111110110101,
	240'b101101101111111111010111010110010101010111001010111111111111111111111111111111111111111111000000010110010101001101010100010101001010110011001000011001011101010111111111111111111111111111111111111111111111111110101011110101011111111110110101,
	240'b101101101111111111010111010110100100111101111110111110001111111111111111111111111111111111111111101100010101010101010100010100110101011110110110110111111110010111111011111111111111111111111111111111111111111111001100110110101111111110110101,
	240'b101101101111111111010111010110100101001101010100101101111111111111111111111111111111111111111111111111011010001101010010010101000101001101011110101011001001010111110101111111111111111111111111111111111111111111100100111000011111111110110101,
	240'b101101101111111111010111010110100101010001010010011001011110000011111111111111111111111111111111111111111111100110010110010100010101010101010100010100000111011011111000111111111111111111111111111111111111111111110011111010001111111110110101,
	240'b101101101111111111010111010110100101010001010101010100010111111011110001111111111111111111111111111111111111111111110100100010100101001101010101010100000111011111111000111111111111111111111111111111111111111111110111111011101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101000010010010111101111111111111111111111111111111111111111111111000010110000001010000010011100111010111111000111111111111111111111111111111111111111111111000111100011111111110110101,
	240'b101101011111111111010111010110100101010001010101010101010101010001010001100101101111011011111111111111111111111111111110101100100110100001101000011001011000011111111001111111111111111111111111111111111111111111111000111100011111111110110101,
	240'b101101011111111111010111010110100101010001010101010101010101010101010100010100101000101111101100111111111111111111111110111100011111000011110000111100001111001111111110111111111111111111111111111111111111111111110100111010101111111110110101,
	240'b101101011111111111010111010110010100111101010000010101000101010101010101010101000101000001110110110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110111001111111110110101,
	240'b101101011111111111010110010111111000001110001010011000100101010001010101010101010101010101010001010111001001100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010001001110101101111111110110101,
	240'b101101011111111111010100011010111110111011111010011111000101000001010101010101010101010101010101010100110101000001100100100101111101000111110011111111111111111111111111111111111111111111111111111100101001011101011010110110101111111110110101,
	240'b101101101111111111010100011010111101100011111111110101000110001101010010010101010101010101010101010101010101010101010011010100000101100101110000100100111010111011000010110011001100110110110011011110000101000101011011110110101111111110110101,
	240'b101101101111111111010110010111111001000011010000111111111100011101011101010101000101010101010101010101010101010101010101010101010101010001010010010100000101000001010101010110000101100001010010010100010101010001011100110110101111111110110101,
	240'b101101101111111111010110010110101100110111001000110101001111111110100111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111010110010110011100010111111110101110101110000011001110010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111010111010101110111011011101011111110001011101010011000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111010111010110100100111110000011111100101111001110111000010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101100111111111111011100010110100101001101010000100101001111111111101010010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110011,
	240'b101001011111110011110101011101100100111001010000011010111011010110100110010101110101000101010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100110101111010111101101111110010100100,
	240'b101011011110010111111111110110000111111101101010011010100110011101100111011010100110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010101000000111011011111111111110001010101100,
	240'b111000001011101111111001111111111111100111110000111100011111000011110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111100111111111111110001011101011100010,
	240'b111100101101010011000000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110101111001101010111110010,
	240'b111110011111110011011101100111001001101010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001100110100001111000111111110011111001,
	240'b111011111111001011101010110000011011000110110011101100111011001010110010101100101011001010110011101100111011001110110011101100111011001110110010101100101011001010110010101100111011001110110011101100111011000110111110111001001111000111101111,
	240'b111100101101111010111101110111111111100111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111100111011101101110001101111011110010,
	240'b111001101011100111110010111111111111111111111010111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110011111100111111001111110101111111111111111111100001011100111101000,
	240'b101100111101111011111111111001111001100101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011111010111110101111101011110010111100101111100011111011001101111101001111111111101110010110010,
	240'b101000111111101011111001100001000100110101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000101010001010100010101000001010111100100111001110101100110010011110100110110000111111110101111101010100001,
	240'b101100101111111111011111010110110101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100001111010111111111010000110010011110101001101011110111000101111111110110001,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101100001110010111111110011100101011100010100111101011100110110101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111100100011100001011111111110110110110011101011010110110101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101110011011101001011000111111111111011100001011001110110101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010010101101111111111111000101110100111101001101011100110110101111111110110101,
	240'b101101101111111111010111010110100101010001010010010100000101001001010010010100000101000001010001010100110101010101010101010101010101010101010101010101010101010101010011011010001101101111111111110000111001001001011111110110101111111110110101,
	240'b101101011111111111010111010110100101000001101001100110101011000010101111101001111001010001111010011000000101001101010001010101000101010101010101010101010101010101010101010100010111001011100100111110101100001101101010110110001111111110110101,
	240'b101101011111111111010111010101111000011111100101111111111111111111111111111111111111111111110111111000011011100010000001010110000101000101010100010101010101010101010101010101010100111110000101111111111110110001101100110110001111111110110101,
	240'b101101011111111111010011011111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011001000000101010100010100100101010101010101010101010101001101101000101000001001010101100011110110011111111110110101,
	240'b101101011111111111010111110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111001011001010101000101010101010101010101010101010100010100010101000001011100110110101111111110110101,
	240'b101101011111111111100111111100111111111111111111111111111111111111111111111111111111101111111010111110101111100111111000111111111111111111111111110111010111100001010001010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111110000111110101111111111111111111111111111111111111111111110011001010101111100011111110111111010111001111111101111111111111111111111111110101110000011010100000101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111110000111110101111111111111111111111111111111111111111111101110111000001001101010011110110001011100100111111111111111111111111111111111111111111101110011111110101000001010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111101101111110011111111111111111111111111111111111111111111101110111001101010001010101010101010010011011111110111111111111111111111111111111111111111111111001100110111101010001010101010101010001011100110110101111111110110101,
	240'b101101101111111111101001111101101111111111111111111111111111111111111111111101110111000101001101010101000101010001010011101010001111111011111111111111111111111111111111111111111100111101011100010100110101010001011100110110101111111110110101,
	240'b101101101111111111100001111001111111111111111111111111111111111111111111111101011000011110010001010101110101010001010011010101111011100011111111111111111111111111111111111111111111111110100101010100010101001101011100110110101111111110110101,
	240'b101101101111111111011000110100101111111111111111111111111111111111111111111110011101110111101010100111110101001001010101010100110101101111000110111111111111111111111111111111111111111111110000011100100101000001011100110110101111111110110101,
	240'b101101011111111111010010101100101111111111111111111111111111111111111111111111111101100101110110110101001001010001010000010101010101001001100010110100111111111111111111111111111111111111111111101111000101001001011100110110101111111110110101,
	240'b101101011111111111010010100011001111110111111111111111111111111111111111111111111010110101001010011101101101100110000110010100000101010101010000011100101110111011111111111111111111111111111111111100110111000001011001110110101111111110110101,
	240'b101101011111111111010101011010001110011011111111111111111111111111111111111111111010000101001111010100001000001011011010011110100101000001010101010100011011111011111111111111111111111111111111111111111010101001011000110110101111111110110101,
	240'b101101011111111111010110010101111011011111111111111111111111111111111111111111111011010001010000010101010101000010010000110110000110111101010001010100001010011011111111111111111111111111111111111111111101110101100101110110011111111110110101,
	240'b101101011111111111010111010101100111101111111001111111111111111111111111111111111110010001100101010100010101010101010001100111101101001101100101010011001010110111111111111111111111111111111111111111111111100110000101110101101111111110110101,
	240'b101101101111111111010111010110010101010111001010111111111111111111111111111111111111111111000000010110010101001101010100010101001010110011001000011001011101010111111111111111111111111111111111111111111111111110101011110101011111111110110101,
	240'b101101101111111111010111010110100100111101111110111110001111111111111111111111111111111111111111101100010101010101010100010100110101011110110110110111111110010111111011111111111111111111111111111111111111111111001100110110101111111110110101,
	240'b101101101111111111010111010110100101001101010100101101111111111111111111111111111111111111111111111111011010001101010010010101000101001101011110101011001001010111110101111111111111111111111111111111111111111111100100111000011111111110110101,
	240'b101101101111111111010111010110100101010001010010011001011110000011111111111111111111111111111111111111111111100110010110010100010101010101010100010100000111011011111000111111111111111111111111111111111111111111110011111010001111111110110101,
	240'b101101101111111111010111010110100101010001010101010100010111111011110001111111111111111111111111111111111111111111110100100010100101001101010101010100000111011111111000111111111111111111111111111111111111111111110111111011101111111110110101,
	240'b101101101111111111010111010110100101010001010101010101010101000010010010111101111111111111111111111111111111111111111111111000010110000001010000010011100111010111111000111111111111111111111111111111111111111111111000111100011111111110110101,
	240'b101101011111111111010111010110100101010001010101010101010101010001010001100101101111011011111111111111111111111111111110101100100110100001101000011001011000011111111001111111111111111111111111111111111111111111111000111100011111111110110101,
	240'b101101011111111111010111010110100101010001010101010101010101010101010100010100101000101111101100111111111111111111111110111100011111000011110000111100001111001111111110111111111111111111111111111111111111111111110100111010101111111110110101,
	240'b101101011111111111010111010110010100111101010000010101000101010101010101010101000101000001110110110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110111001111111110110101,
	240'b101101011111111111010110010111111000001110001010011000100101010001010101010101010101010101010001010111001001100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010001001110101101111111110110101,
	240'b101101011111111111010100011010111110111011111010011111000101000001010101010101010101010101010101010100110101000001100100100101111101000111110011111111111111111111111111111111111111111111111111111100101001011101011010110110101111111110110101,
	240'b101101101111111111010100011010111101100011111111110101000110001101010010010101010101010101010101010101010101010101010011010100000101100101110000100100111010111011000010110011001100110110110011011110000101000101011011110110101111111110110101,
	240'b101101101111111111010110010111111001000011010000111111111100011101011101010101000101010101010101010101010101010101010101010101010101010001010010010100000101000001010101010110000101100001010010010100010101010001011100110110101111111110110101,
	240'b101101101111111111010110010110101100110111001000110101001111111110100111010100010101010101010101010101010101010101010101010101010101010101010101010101010101010101010100010101000101010001010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111010110010110011100010111111110101110101110000011001110010101100101010001010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111010111010101110111011011101011111110001011101010011000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101101101111111111010111010110100100111110000011111100101111001110111000010111010101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001011100110110101111111110110101,
	240'b101100111111111111011100010110100101001101010000100101001111111111101010010111100101001101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101001101011101110111111111111110110011,
	240'b101001011111110011110101011101100100111001010000011010111011010110100110010101110101000101010010010100100101001001010010010100100101001001010010010100100101001001010010010100100101001001010010010100100100110101111010111101101111110010100100,
	240'b101011011110010111111111110110000111111101101010011010100110011101100111011010100110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010110110101101101011011010101000000111011011111111111110001010101100,
	240'b111000001011101111111001111111111111100111110000111100011111000011110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111000111110001111100011111100111111111111110001011101011100010,
	240'b111100101101010011000000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110101111001101010111110010,
	240'b111110011111110011011101100111001001101010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101100001011000010110000101011111001100110100001111000111111110011111001,
};
always_comb begin
	if((x_pin <= x_cnt && x_cnt <= x_pin + X_WIDTH) && (y_pin <= y_cnt && y_cnt <= y_pin + Y_WIDTH)) begin
		r_data = picture[(y_cnt - y_pin)][(x_cnt - x_pin)<<3 +: 8];
		g_data = picture[(y_cnt - y_pin) + Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
		b_data = picture[(y_cnt - y_pin) + 2*Y_WIDTH][(x_cnt - x_pin)<<3 +: 8];
	end
	else begin
		r_data = 8'b0;
		g_data = 8'b0;
		b_data = 8'b0;
	end
end
endmodule